-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d3",
     9 => x"a4080b0b",
    10 => x"80d3a808",
    11 => x"0b0b80d3",
    12 => x"ac080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d3ac0c0b",
    16 => x"0b80d3a8",
    17 => x"0c0b0b80",
    18 => x"d3a40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbdd0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d3a470",
    57 => x"80dde427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518a8f",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d3",
    65 => x"b40c9f0b",
    66 => x"80d3b80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d3b808ff",
    70 => x"0580d3b8",
    71 => x"0c80d3b8",
    72 => x"088025e8",
    73 => x"3880d3b4",
    74 => x"08ff0580",
    75 => x"d3b40c80",
    76 => x"d3b40880",
    77 => x"25d03880",
    78 => x"0b80d3b8",
    79 => x"0c800b80",
    80 => x"d3b40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d3b408",
   100 => x"25913882",
   101 => x"c82d80d3",
   102 => x"b408ff05",
   103 => x"80d3b40c",
   104 => x"838a0480",
   105 => x"d3b40880",
   106 => x"d3b80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d3b408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d3b80881",
   116 => x"0580d3b8",
   117 => x"0c80d3b8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d3b8",
   121 => x"0c80d3b4",
   122 => x"08810580",
   123 => x"d3b40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d3",
   128 => x"b8088105",
   129 => x"80d3b80c",
   130 => x"80d3b808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d3b8",
   134 => x"0c80d3b4",
   135 => x"08810580",
   136 => x"d3b40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d3bc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d3bc0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d3",
   177 => x"bc088407",
   178 => x"80d3bc0c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5483f474",
   182 => x"258f3883",
   183 => x"0b0b0b80",
   184 => x"cab80c82",
   185 => x"845385f3",
   186 => x"04810b0b",
   187 => x"0b80cab8",
   188 => x"0ca8530b",
   189 => x"0b80cab8",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0c747431",
   193 => x"ffb005ff",
   194 => x"1271712c",
   195 => x"ff941970",
   196 => x"9f2a1170",
   197 => x"812c80d3",
   198 => x"bc085255",
   199 => x"51525652",
   200 => x"53517680",
   201 => x"2e853870",
   202 => x"81075170",
   203 => x"f6940c72",
   204 => x"098105f6",
   205 => x"800c7109",
   206 => x"8105f684",
   207 => x"0c029405",
   208 => x"0d040402",
   209 => x"fc050d80",
   210 => x"cfc85194",
   211 => x"b52d0284",
   212 => x"050d0402",
   213 => x"fc050d80",
   214 => x"cabc5194",
   215 => x"b52d0284",
   216 => x"050d0402",
   217 => x"fc050d80",
   218 => x"cea05194",
   219 => x"b52d0284",
   220 => x"050d0402",
   221 => x"fc050d81",
   222 => x"808051c0",
   223 => x"115170fb",
   224 => x"38028405",
   225 => x"0d047181",
   226 => x"2e098106",
   227 => x"893881c3",
   228 => x"0bec0c87",
   229 => x"9a04830b",
   230 => x"ec0c86f3",
   231 => x"2d820bec",
   232 => x"0c0491fd",
   233 => x"2d80d3a4",
   234 => x"0880ce90",
   235 => x"0c91fd2d",
   236 => x"80d3a408",
   237 => x"80cdbc0c",
   238 => x"91fd2d80",
   239 => x"d3a40880",
   240 => x"d0e00c91",
   241 => x"fd2d80d3",
   242 => x"a40880cf",
   243 => x"b80c91fd",
   244 => x"2d80d3a4",
   245 => x"0880cbe0",
   246 => x"0c0402fc",
   247 => x"050d84bf",
   248 => x"5186f32d",
   249 => x"ff115170",
   250 => x"8025f638",
   251 => x"0284050d",
   252 => x"0402f405",
   253 => x"0d745372",
   254 => x"70810554",
   255 => x"80f52d52",
   256 => x"71802e89",
   257 => x"38715183",
   258 => x"842d87f7",
   259 => x"04810b80",
   260 => x"d3a40c02",
   261 => x"8c050d04",
   262 => x"02dc050d",
   263 => x"80598184",
   264 => x"0bec0c7a",
   265 => x"5280d3c0",
   266 => x"51b38d2d",
   267 => x"80d3a408",
   268 => x"792e819b",
   269 => x"3880d3c4",
   270 => x"08547385",
   271 => x"2e098106",
   272 => x"8a38840b",
   273 => x"ec0c8153",
   274 => x"89d70473",
   275 => x"f80c81a4",
   276 => x"0bec0c87",
   277 => x"da2d78ff",
   278 => x"15565874",
   279 => x"802e8b38",
   280 => x"81187581",
   281 => x"2a565888",
   282 => x"db04f718",
   283 => x"58815980",
   284 => x"742580d7",
   285 => x"38a40bec",
   286 => x"0c775274",
   287 => x"5184a82d",
   288 => x"80d49c52",
   289 => x"80d3c051",
   290 => x"b6802d80",
   291 => x"d3a40880",
   292 => x"2ea03880",
   293 => x"d49c5783",
   294 => x"fc567670",
   295 => x"84055808",
   296 => x"e80cfc16",
   297 => x"56758025",
   298 => x"f13881a4",
   299 => x"0bec0c89",
   300 => x"ba0480d3",
   301 => x"a4085984",
   302 => x"805480d3",
   303 => x"c051b5d0",
   304 => x"2dfc8014",
   305 => x"81165654",
   306 => x"88ef0484",
   307 => x"0bec0c80",
   308 => x"d3c408f8",
   309 => x"0c785372",
   310 => x"80d3a40c",
   311 => x"02a4050d",
   312 => x"0402f805",
   313 => x"0d735188",
   314 => x"982d80d3",
   315 => x"a4085280",
   316 => x"d3a40880",
   317 => x"2e883880",
   318 => x"cdcc518a",
   319 => x"820480cd",
   320 => x"a85194b5",
   321 => x"2d7180d3",
   322 => x"a40c0288",
   323 => x"050d0402",
   324 => x"f0050d80",
   325 => x"0b80d3cc",
   326 => x"0c815187",
   327 => x"862d8051",
   328 => x"87862d84",
   329 => x"0bec0c91",
   330 => x"cd2d8df8",
   331 => x"2d81f92d",
   332 => x"835291b0",
   333 => x"2d815185",
   334 => x"8d2dff12",
   335 => x"52718025",
   336 => x"f13880c4",
   337 => x"0bec0c80",
   338 => x"c8985187",
   339 => x"f12da9c5",
   340 => x"2d80d3a4",
   341 => x"08802e83",
   342 => x"88388184",
   343 => x"0bec0c80",
   344 => x"c8b05187",
   345 => x"f12d80d3",
   346 => x"cc08bfff",
   347 => x"ff068780",
   348 => x"077080d3",
   349 => x"cc0cfc0c",
   350 => x"80c8c851",
   351 => x"88982d80",
   352 => x"d3a40880",
   353 => x"2eac3880",
   354 => x"c8d45188",
   355 => x"982d80d3",
   356 => x"a408802e",
   357 => x"9d3880c8",
   358 => x"e0518898",
   359 => x"2d80d3a4",
   360 => x"08802e8e",
   361 => x"38805187",
   362 => x"862d8051",
   363 => x"858d2d8b",
   364 => x"b90480c8",
   365 => x"ec5187f1",
   366 => x"2d840bec",
   367 => x"0c89e151",
   368 => x"bdca2d80",
   369 => x"d3cc0880",
   370 => x"d1b80c80",
   371 => x"d3cc08fc",
   372 => x"0c80ccb0",
   373 => x"0b80d3d0",
   374 => x"0c80ccb0",
   375 => x"5194b52d",
   376 => x"805187a2",
   377 => x"2d830b80",
   378 => x"d4900c92",
   379 => x"862d8051",
   380 => x"858d2d92",
   381 => x"9a2d8e84",
   382 => x"2d94c82d",
   383 => x"80cadc0b",
   384 => x"80f52d80",
   385 => x"cae80b80",
   386 => x"f52d718a",
   387 => x"2b718b2b",
   388 => x"0780cb80",
   389 => x"0b80f52d",
   390 => x"708d2b72",
   391 => x"0780cb98",
   392 => x"0b80f52d",
   393 => x"708e2b72",
   394 => x"0780cbc8",
   395 => x"0b80f52d",
   396 => x"70912b72",
   397 => x"077080d3",
   398 => x"cc0c80d1",
   399 => x"b8087081",
   400 => x"06545253",
   401 => x"54525452",
   402 => x"53545553",
   403 => x"71802e88",
   404 => x"38738107",
   405 => x"80d3cc0c",
   406 => x"72812a70",
   407 => x"81065152",
   408 => x"71802e8b",
   409 => x"3880d3cc",
   410 => x"08820780",
   411 => x"d3cc0c72",
   412 => x"822a7081",
   413 => x"06515271",
   414 => x"802e8b38",
   415 => x"80d3cc08",
   416 => x"840780d3",
   417 => x"cc0c7283",
   418 => x"2a708106",
   419 => x"51527180",
   420 => x"2e8b3880",
   421 => x"d3cc0888",
   422 => x"0780d3cc",
   423 => x"0c72842a",
   424 => x"70810651",
   425 => x"5271802e",
   426 => x"8b3880d3",
   427 => x"cc089007",
   428 => x"80d3cc0c",
   429 => x"72852a70",
   430 => x"81065152",
   431 => x"71802e8b",
   432 => x"3880d3cc",
   433 => x"08a00780",
   434 => x"d3cc0c80",
   435 => x"d3cc08fc",
   436 => x"0c865280",
   437 => x"d3a40883",
   438 => x"38845271",
   439 => x"ec0c8bf6",
   440 => x"04800b80",
   441 => x"d3a40c02",
   442 => x"90050d04",
   443 => x"71980c04",
   444 => x"ffb00880",
   445 => x"d3a40c04",
   446 => x"810bffb0",
   447 => x"0c04800b",
   448 => x"ffb00c04",
   449 => x"02f4050d",
   450 => x"8f920480",
   451 => x"d3a40881",
   452 => x"f02e0981",
   453 => x"068a3881",
   454 => x"0b80d1b0",
   455 => x"0c8f9204",
   456 => x"80d3a408",
   457 => x"81e02e09",
   458 => x"81068a38",
   459 => x"810b80d1",
   460 => x"b40c8f92",
   461 => x"0480d3a4",
   462 => x"085280d1",
   463 => x"b408802e",
   464 => x"893880d3",
   465 => x"a4088180",
   466 => x"05527184",
   467 => x"2c728f06",
   468 => x"535380d1",
   469 => x"b008802e",
   470 => x"9a387284",
   471 => x"2980d0f0",
   472 => x"05721381",
   473 => x"712b7009",
   474 => x"73080673",
   475 => x"0c515353",
   476 => x"8f860472",
   477 => x"842980d0",
   478 => x"f0057213",
   479 => x"83712b72",
   480 => x"0807720c",
   481 => x"5353800b",
   482 => x"80d1b40c",
   483 => x"800b80d1",
   484 => x"b00c80d3",
   485 => x"d4519099",
   486 => x"2d80d3a4",
   487 => x"08ff24fe",
   488 => x"ea38800b",
   489 => x"80d3a40c",
   490 => x"028c050d",
   491 => x"0402f805",
   492 => x"0d80d0f0",
   493 => x"528f5180",
   494 => x"72708405",
   495 => x"540cff11",
   496 => x"51708025",
   497 => x"f2380288",
   498 => x"050d0402",
   499 => x"f0050d75",
   500 => x"518dfe2d",
   501 => x"70822cfc",
   502 => x"0680d0f0",
   503 => x"1172109e",
   504 => x"06710870",
   505 => x"722a7083",
   506 => x"0682742b",
   507 => x"70097406",
   508 => x"760c5451",
   509 => x"56575351",
   510 => x"538df82d",
   511 => x"7180d3a4",
   512 => x"0c029005",
   513 => x"0d0402fc",
   514 => x"050d7251",
   515 => x"80710c80",
   516 => x"0b84120c",
   517 => x"0284050d",
   518 => x"0402f005",
   519 => x"0d757008",
   520 => x"84120853",
   521 => x"5353ff54",
   522 => x"71712ea8",
   523 => x"388dfe2d",
   524 => x"84130870",
   525 => x"84291488",
   526 => x"11700870",
   527 => x"81ff0684",
   528 => x"18088111",
   529 => x"8706841a",
   530 => x"0c535155",
   531 => x"5151518d",
   532 => x"f82d7154",
   533 => x"7380d3a4",
   534 => x"0c029005",
   535 => x"0d0402f4",
   536 => x"050d8dfe",
   537 => x"2de00870",
   538 => x"8b2a7081",
   539 => x"06515253",
   540 => x"70802ea1",
   541 => x"3880d3d4",
   542 => x"08708429",
   543 => x"80d3dc05",
   544 => x"7481ff06",
   545 => x"710c5151",
   546 => x"80d3d408",
   547 => x"81118706",
   548 => x"80d3d40c",
   549 => x"51728c2c",
   550 => x"83ff0680",
   551 => x"d3fc0c80",
   552 => x"0b80d480",
   553 => x"0c8df02d",
   554 => x"8df82d02",
   555 => x"8c050d04",
   556 => x"02fc050d",
   557 => x"8dfe2d81",
   558 => x"0b80d480",
   559 => x"0c8df82d",
   560 => x"80d48008",
   561 => x"5170f938",
   562 => x"0284050d",
   563 => x"0402fc05",
   564 => x"0d80d3d4",
   565 => x"5190862d",
   566 => x"8fad2d90",
   567 => x"de518dec",
   568 => x"2d028405",
   569 => x"0d0402fc",
   570 => x"050d8fcf",
   571 => x"5186f32d",
   572 => x"ff115170",
   573 => x"8025f638",
   574 => x"0284050d",
   575 => x"0480d488",
   576 => x"0880d3a4",
   577 => x"0c0402fc",
   578 => x"050d810b",
   579 => x"80d1e40c",
   580 => x"8151858d",
   581 => x"2d028405",
   582 => x"0d0402fc",
   583 => x"050d92a4",
   584 => x"048e842d",
   585 => x"80f6518f",
   586 => x"cb2d80d3",
   587 => x"a408f238",
   588 => x"80da518f",
   589 => x"cb2d80d3",
   590 => x"a408e638",
   591 => x"80d1e008",
   592 => x"518fcb2d",
   593 => x"80d3a408",
   594 => x"d83880d3",
   595 => x"a40880d1",
   596 => x"e40c80d3",
   597 => x"a4085185",
   598 => x"8d2d0284",
   599 => x"050d0402",
   600 => x"ec050d76",
   601 => x"54805287",
   602 => x"0b881580",
   603 => x"f52d5653",
   604 => x"74722483",
   605 => x"38a05372",
   606 => x"5183842d",
   607 => x"81128b15",
   608 => x"80f52d54",
   609 => x"52727225",
   610 => x"de380294",
   611 => x"050d0402",
   612 => x"f0050d80",
   613 => x"d4880854",
   614 => x"81f92d80",
   615 => x"0b80d48c",
   616 => x"0c730880",
   617 => x"2e818938",
   618 => x"820b80d3",
   619 => x"b80c80d4",
   620 => x"8c088f06",
   621 => x"80d3b40c",
   622 => x"73085271",
   623 => x"832e9638",
   624 => x"71832689",
   625 => x"3871812e",
   626 => x"b0389499",
   627 => x"0471852e",
   628 => x"a0389499",
   629 => x"04881480",
   630 => x"f52d8415",
   631 => x"0880c984",
   632 => x"53545287",
   633 => x"f12d7184",
   634 => x"29137008",
   635 => x"5252949d",
   636 => x"04735192",
   637 => x"df2d9499",
   638 => x"0480d1b8",
   639 => x"08881508",
   640 => x"2c708106",
   641 => x"51527180",
   642 => x"2e883880",
   643 => x"c9885194",
   644 => x"960480c9",
   645 => x"8c5187f1",
   646 => x"2d841408",
   647 => x"5187f12d",
   648 => x"80d48c08",
   649 => x"810580d4",
   650 => x"8c0c8c14",
   651 => x"5493a104",
   652 => x"0290050d",
   653 => x"047180d4",
   654 => x"880c938f",
   655 => x"2d80d48c",
   656 => x"08ff0580",
   657 => x"d4900c04",
   658 => x"02e8050d",
   659 => x"80d48808",
   660 => x"80d49408",
   661 => x"575580f6",
   662 => x"518fcb2d",
   663 => x"80d3a408",
   664 => x"812a7081",
   665 => x"06515271",
   666 => x"802ea238",
   667 => x"94f2048e",
   668 => x"842d80f6",
   669 => x"518fcb2d",
   670 => x"80d3a408",
   671 => x"f23880d1",
   672 => x"e4088132",
   673 => x"7080d1e4",
   674 => x"0c51858d",
   675 => x"2d800b80",
   676 => x"d4840c8c",
   677 => x"518fcb2d",
   678 => x"80d3a408",
   679 => x"812a7081",
   680 => x"06515271",
   681 => x"802e80d1",
   682 => x"3880d1bc",
   683 => x"0880d1d0",
   684 => x"0880d1bc",
   685 => x"0c80d1d0",
   686 => x"0c80d1c0",
   687 => x"0880d1d4",
   688 => x"0880d1c0",
   689 => x"0c80d1d4",
   690 => x"0c80d1c4",
   691 => x"0880d1d8",
   692 => x"0880d1c4",
   693 => x"0c80d1d8",
   694 => x"0c80d1c8",
   695 => x"0880d1dc",
   696 => x"0880d1c8",
   697 => x"0c80d1dc",
   698 => x"0c80d1cc",
   699 => x"0880d1e0",
   700 => x"0880d1cc",
   701 => x"0c80d1e0",
   702 => x"0c80d3fc",
   703 => x"08a00652",
   704 => x"80722596",
   705 => x"3891e62d",
   706 => x"8e842d80",
   707 => x"d1e40881",
   708 => x"327080d1",
   709 => x"e40c5185",
   710 => x"8d2d80d1",
   711 => x"e40882ef",
   712 => x"3880d1d0",
   713 => x"08518fcb",
   714 => x"2d80d3a4",
   715 => x"08802e8b",
   716 => x"3880d484",
   717 => x"08810780",
   718 => x"d4840c80",
   719 => x"d1d40851",
   720 => x"8fcb2d80",
   721 => x"d3a40880",
   722 => x"2e8b3880",
   723 => x"d4840882",
   724 => x"0780d484",
   725 => x"0c80d1d8",
   726 => x"08518fcb",
   727 => x"2d80d3a4",
   728 => x"08802e8b",
   729 => x"3880d484",
   730 => x"08840780",
   731 => x"d4840c80",
   732 => x"d1dc0851",
   733 => x"8fcb2d80",
   734 => x"d3a40880",
   735 => x"2e8b3880",
   736 => x"d4840888",
   737 => x"0780d484",
   738 => x"0c80d1e0",
   739 => x"08518fcb",
   740 => x"2d80d3a4",
   741 => x"08802e8b",
   742 => x"3880d484",
   743 => x"08900780",
   744 => x"d4840c80",
   745 => x"d1bc0851",
   746 => x"8fcb2d80",
   747 => x"d3a40880",
   748 => x"2e8c3880",
   749 => x"d4840882",
   750 => x"800780d4",
   751 => x"840c80d1",
   752 => x"c008518f",
   753 => x"cb2d80d3",
   754 => x"a408802e",
   755 => x"8c3880d4",
   756 => x"84088480",
   757 => x"0780d484",
   758 => x"0c80d1c4",
   759 => x"08518fcb",
   760 => x"2d80d3a4",
   761 => x"08802e8c",
   762 => x"3880d484",
   763 => x"08888007",
   764 => x"80d4840c",
   765 => x"80d1c808",
   766 => x"518fcb2d",
   767 => x"80d3a408",
   768 => x"802e8c38",
   769 => x"80d48408",
   770 => x"90800780",
   771 => x"d4840c80",
   772 => x"d1cc0851",
   773 => x"8fcb2d80",
   774 => x"d3a40880",
   775 => x"2e8c3880",
   776 => x"d48408a0",
   777 => x"800780d4",
   778 => x"840c9451",
   779 => x"8fcb2d80",
   780 => x"d3a40852",
   781 => x"91518fcb",
   782 => x"2d7180d3",
   783 => x"a4080652",
   784 => x"80e6518f",
   785 => x"cb2d7180",
   786 => x"d3a40806",
   787 => x"5271802e",
   788 => x"8d3880d4",
   789 => x"84088480",
   790 => x"800780d4",
   791 => x"840c80fe",
   792 => x"518fcb2d",
   793 => x"80d3a408",
   794 => x"5287518f",
   795 => x"cb2d7180",
   796 => x"d3a40807",
   797 => x"5271802e",
   798 => x"8d3880d4",
   799 => x"84088880",
   800 => x"800780d4",
   801 => x"840c80d4",
   802 => x"8408ed0c",
   803 => x"a19a0494",
   804 => x"518fcb2d",
   805 => x"80d3a408",
   806 => x"5291518f",
   807 => x"cb2d7180",
   808 => x"d3a40806",
   809 => x"5280e651",
   810 => x"8fcb2d71",
   811 => x"80d3a408",
   812 => x"06527180",
   813 => x"2e8d3880",
   814 => x"d4840884",
   815 => x"80800780",
   816 => x"d4840c80",
   817 => x"fe518fcb",
   818 => x"2d80d3a4",
   819 => x"08528751",
   820 => x"8fcb2d71",
   821 => x"80d3a408",
   822 => x"07527180",
   823 => x"2e8d3880",
   824 => x"d4840888",
   825 => x"80800780",
   826 => x"d4840c80",
   827 => x"d48408ed",
   828 => x"0c81f551",
   829 => x"8fcb2d80",
   830 => x"d3a40881",
   831 => x"2a708106",
   832 => x"515271a4",
   833 => x"3880d1d0",
   834 => x"08518fcb",
   835 => x"2d80d3a4",
   836 => x"08812a70",
   837 => x"81065152",
   838 => x"718e3880",
   839 => x"d3fc0881",
   840 => x"06528072",
   841 => x"2580c238",
   842 => x"80d3fc08",
   843 => x"81065280",
   844 => x"72258438",
   845 => x"91e62d80",
   846 => x"d4900852",
   847 => x"71802e8a",
   848 => x"38ff1280",
   849 => x"d4900c9a",
   850 => x"e90480d4",
   851 => x"8c081080",
   852 => x"d48c0805",
   853 => x"70842916",
   854 => x"51528812",
   855 => x"08802e89",
   856 => x"38ff5188",
   857 => x"12085271",
   858 => x"2d81f251",
   859 => x"8fcb2d80",
   860 => x"d3a40881",
   861 => x"2a708106",
   862 => x"515271a4",
   863 => x"3880d1d4",
   864 => x"08518fcb",
   865 => x"2d80d3a4",
   866 => x"08812a70",
   867 => x"81065152",
   868 => x"718e3880",
   869 => x"d3fc0882",
   870 => x"06528072",
   871 => x"2580c338",
   872 => x"80d3fc08",
   873 => x"82065280",
   874 => x"72258438",
   875 => x"91e62d80",
   876 => x"d48c08ff",
   877 => x"1180d490",
   878 => x"08565353",
   879 => x"7372258a",
   880 => x"38811480",
   881 => x"d4900c9b",
   882 => x"e2047210",
   883 => x"13708429",
   884 => x"16515288",
   885 => x"1208802e",
   886 => x"8938fe51",
   887 => x"88120852",
   888 => x"712d81fd",
   889 => x"518fcb2d",
   890 => x"80d3a408",
   891 => x"812a7081",
   892 => x"06515271",
   893 => x"a43880d1",
   894 => x"d808518f",
   895 => x"cb2d80d3",
   896 => x"a408812a",
   897 => x"70810651",
   898 => x"52718e38",
   899 => x"80d3fc08",
   900 => x"84065280",
   901 => x"722580c0",
   902 => x"3880d3fc",
   903 => x"08840652",
   904 => x"80722584",
   905 => x"3891e62d",
   906 => x"80d49008",
   907 => x"802e8a38",
   908 => x"800b80d4",
   909 => x"900c9cd8",
   910 => x"0480d48c",
   911 => x"081080d4",
   912 => x"8c080570",
   913 => x"84291651",
   914 => x"52881208",
   915 => x"802e8938",
   916 => x"fd518812",
   917 => x"0852712d",
   918 => x"81fa518f",
   919 => x"cb2d80d3",
   920 => x"a408812a",
   921 => x"70810651",
   922 => x"5271a438",
   923 => x"80d1dc08",
   924 => x"518fcb2d",
   925 => x"80d3a408",
   926 => x"812a7081",
   927 => x"06515271",
   928 => x"8e3880d3",
   929 => x"fc088806",
   930 => x"52807225",
   931 => x"80c03880",
   932 => x"d3fc0888",
   933 => x"06528072",
   934 => x"25843891",
   935 => x"e62d80d4",
   936 => x"8c08ff11",
   937 => x"545280d4",
   938 => x"90087325",
   939 => x"89387280",
   940 => x"d4900c9d",
   941 => x"ce047110",
   942 => x"12708429",
   943 => x"16515288",
   944 => x"1208802e",
   945 => x"8938fc51",
   946 => x"88120852",
   947 => x"712d80d4",
   948 => x"90087053",
   949 => x"5473802e",
   950 => x"8a388c15",
   951 => x"ff155555",
   952 => x"9dd50482",
   953 => x"0b80d3b8",
   954 => x"0c718f06",
   955 => x"80d3b40c",
   956 => x"81eb518f",
   957 => x"cb2d80d3",
   958 => x"a408812a",
   959 => x"70810651",
   960 => x"5271802e",
   961 => x"ad387408",
   962 => x"852e0981",
   963 => x"06a43888",
   964 => x"1580f52d",
   965 => x"ff055271",
   966 => x"881681b7",
   967 => x"2d71982b",
   968 => x"52718025",
   969 => x"8838800b",
   970 => x"881681b7",
   971 => x"2d745192",
   972 => x"df2d81f4",
   973 => x"518fcb2d",
   974 => x"80d3a408",
   975 => x"812a7081",
   976 => x"06515271",
   977 => x"802eb338",
   978 => x"7408852e",
   979 => x"098106aa",
   980 => x"38881580",
   981 => x"f52d8105",
   982 => x"52718816",
   983 => x"81b72d71",
   984 => x"81ff068b",
   985 => x"1680f52d",
   986 => x"54527272",
   987 => x"27873872",
   988 => x"881681b7",
   989 => x"2d745192",
   990 => x"df2d80da",
   991 => x"518fcb2d",
   992 => x"80d3a408",
   993 => x"812a7081",
   994 => x"06515271",
   995 => x"8e3880d3",
   996 => x"fc089006",
   997 => x"52807225",
   998 => x"81bc3880",
   999 => x"d4880880",
  1000 => x"d3fc0890",
  1001 => x"06535380",
  1002 => x"72258438",
  1003 => x"91e62d80",
  1004 => x"d4900854",
  1005 => x"73802e8a",
  1006 => x"388c13ff",
  1007 => x"1555539f",
  1008 => x"b4047208",
  1009 => x"5271822e",
  1010 => x"a6387182",
  1011 => x"26893871",
  1012 => x"812eaa38",
  1013 => x"a0d60471",
  1014 => x"832eb438",
  1015 => x"71842e09",
  1016 => x"810680f2",
  1017 => x"38881308",
  1018 => x"5194b52d",
  1019 => x"a0d60480",
  1020 => x"d4900851",
  1021 => x"88130852",
  1022 => x"712da0d6",
  1023 => x"04810b88",
  1024 => x"14082b80",
  1025 => x"d1b80832",
  1026 => x"80d1b80c",
  1027 => x"a0aa0488",
  1028 => x"1380f52d",
  1029 => x"81058b14",
  1030 => x"80f52d53",
  1031 => x"54717424",
  1032 => x"83388054",
  1033 => x"73881481",
  1034 => x"b72d938f",
  1035 => x"2da0d604",
  1036 => x"7508802e",
  1037 => x"a4387508",
  1038 => x"518fcb2d",
  1039 => x"80d3a408",
  1040 => x"81065271",
  1041 => x"802e8c38",
  1042 => x"80d49008",
  1043 => x"51841608",
  1044 => x"52712d88",
  1045 => x"165675d8",
  1046 => x"38805480",
  1047 => x"0b80d3b8",
  1048 => x"0c738f06",
  1049 => x"80d3b40c",
  1050 => x"a0527380",
  1051 => x"d490082e",
  1052 => x"09810699",
  1053 => x"3880d48c",
  1054 => x"08ff0574",
  1055 => x"32700981",
  1056 => x"05707207",
  1057 => x"9f2a9171",
  1058 => x"31515153",
  1059 => x"53715183",
  1060 => x"842d8114",
  1061 => x"548e7425",
  1062 => x"c23880d1",
  1063 => x"e40880d3",
  1064 => x"a40c0298",
  1065 => x"050d0402",
  1066 => x"f4050dd4",
  1067 => x"5281ff72",
  1068 => x"0c710853",
  1069 => x"81ff720c",
  1070 => x"72882b83",
  1071 => x"fe800672",
  1072 => x"087081ff",
  1073 => x"06515253",
  1074 => x"81ff720c",
  1075 => x"72710788",
  1076 => x"2b720870",
  1077 => x"81ff0651",
  1078 => x"525381ff",
  1079 => x"720c7271",
  1080 => x"07882b72",
  1081 => x"087081ff",
  1082 => x"06720780",
  1083 => x"d3a40c52",
  1084 => x"53028c05",
  1085 => x"0d0402f4",
  1086 => x"050d7476",
  1087 => x"7181ff06",
  1088 => x"d40c5353",
  1089 => x"80d49808",
  1090 => x"85387189",
  1091 => x"2b527198",
  1092 => x"2ad40c71",
  1093 => x"902a7081",
  1094 => x"ff06d40c",
  1095 => x"5171882a",
  1096 => x"7081ff06",
  1097 => x"d40c5171",
  1098 => x"81ff06d4",
  1099 => x"0c72902a",
  1100 => x"7081ff06",
  1101 => x"d40c51d4",
  1102 => x"087081ff",
  1103 => x"06515182",
  1104 => x"b8bf5270",
  1105 => x"81ff2e09",
  1106 => x"81069438",
  1107 => x"81ff0bd4",
  1108 => x"0cd40870",
  1109 => x"81ff06ff",
  1110 => x"14545151",
  1111 => x"71e53870",
  1112 => x"80d3a40c",
  1113 => x"028c050d",
  1114 => x"0402fc05",
  1115 => x"0d81c751",
  1116 => x"81ff0bd4",
  1117 => x"0cff1151",
  1118 => x"708025f4",
  1119 => x"38028405",
  1120 => x"0d0402f4",
  1121 => x"050d81ff",
  1122 => x"0bd40c93",
  1123 => x"53805287",
  1124 => x"fc80c151",
  1125 => x"a1f62d80",
  1126 => x"d3a4088b",
  1127 => x"3881ff0b",
  1128 => x"d40c8153",
  1129 => x"a3b004a2",
  1130 => x"e92dff13",
  1131 => x"5372de38",
  1132 => x"7280d3a4",
  1133 => x"0c028c05",
  1134 => x"0d0402ec",
  1135 => x"050d810b",
  1136 => x"80d4980c",
  1137 => x"8454d008",
  1138 => x"708f2a70",
  1139 => x"81065151",
  1140 => x"5372f338",
  1141 => x"72d00ca2",
  1142 => x"e92d80c9",
  1143 => x"905187f1",
  1144 => x"2dd00870",
  1145 => x"8f2a7081",
  1146 => x"06515153",
  1147 => x"72f33881",
  1148 => x"0bd00cb1",
  1149 => x"53805284",
  1150 => x"d480c051",
  1151 => x"a1f62d80",
  1152 => x"d3a40881",
  1153 => x"2e933872",
  1154 => x"822ebf38",
  1155 => x"ff135372",
  1156 => x"e438ff14",
  1157 => x"5473ffae",
  1158 => x"38a2e92d",
  1159 => x"83aa5284",
  1160 => x"9c80c851",
  1161 => x"a1f62d80",
  1162 => x"d3a40881",
  1163 => x"2e098106",
  1164 => x"9338a1a7",
  1165 => x"2d80d3a4",
  1166 => x"0883ffff",
  1167 => x"06537283",
  1168 => x"aa2e9f38",
  1169 => x"a3822da4",
  1170 => x"dd0480c9",
  1171 => x"9c5187f1",
  1172 => x"2d8053a6",
  1173 => x"b20480c9",
  1174 => x"b45187f1",
  1175 => x"2d8054a6",
  1176 => x"830481ff",
  1177 => x"0bd40cb1",
  1178 => x"54a2e92d",
  1179 => x"8fcf5380",
  1180 => x"5287fc80",
  1181 => x"f751a1f6",
  1182 => x"2d80d3a4",
  1183 => x"085580d3",
  1184 => x"a408812e",
  1185 => x"0981069c",
  1186 => x"3881ff0b",
  1187 => x"d40c820a",
  1188 => x"52849c80",
  1189 => x"e951a1f6",
  1190 => x"2d80d3a4",
  1191 => x"08802e8d",
  1192 => x"38a2e92d",
  1193 => x"ff135372",
  1194 => x"c638a5f6",
  1195 => x"0481ff0b",
  1196 => x"d40c80d3",
  1197 => x"a4085287",
  1198 => x"fc80fa51",
  1199 => x"a1f62d80",
  1200 => x"d3a408b2",
  1201 => x"3881ff0b",
  1202 => x"d40cd408",
  1203 => x"5381ff0b",
  1204 => x"d40c81ff",
  1205 => x"0bd40c81",
  1206 => x"ff0bd40c",
  1207 => x"81ff0bd4",
  1208 => x"0c72862a",
  1209 => x"70810676",
  1210 => x"56515372",
  1211 => x"963880d3",
  1212 => x"a40854a6",
  1213 => x"83047382",
  1214 => x"2efedb38",
  1215 => x"ff145473",
  1216 => x"fee73873",
  1217 => x"80d4980c",
  1218 => x"738b3881",
  1219 => x"5287fc80",
  1220 => x"d051a1f6",
  1221 => x"2d81ff0b",
  1222 => x"d40cd008",
  1223 => x"708f2a70",
  1224 => x"81065151",
  1225 => x"5372f338",
  1226 => x"72d00c81",
  1227 => x"ff0bd40c",
  1228 => x"81537280",
  1229 => x"d3a40c02",
  1230 => x"94050d04",
  1231 => x"02e8050d",
  1232 => x"78558056",
  1233 => x"81ff0bd4",
  1234 => x"0cd00870",
  1235 => x"8f2a7081",
  1236 => x"06515153",
  1237 => x"72f33882",
  1238 => x"810bd00c",
  1239 => x"81ff0bd4",
  1240 => x"0c775287",
  1241 => x"fc80d151",
  1242 => x"a1f62d80",
  1243 => x"dbc6df54",
  1244 => x"80d3a408",
  1245 => x"802e8b38",
  1246 => x"80c9d451",
  1247 => x"87f12da7",
  1248 => x"d60481ff",
  1249 => x"0bd40cd4",
  1250 => x"087081ff",
  1251 => x"06515372",
  1252 => x"81fe2e09",
  1253 => x"81069e38",
  1254 => x"80ff53a1",
  1255 => x"a72d80d3",
  1256 => x"a4087570",
  1257 => x"8405570c",
  1258 => x"ff135372",
  1259 => x"8025ec38",
  1260 => x"8156a7bb",
  1261 => x"04ff1454",
  1262 => x"73c83881",
  1263 => x"ff0bd40c",
  1264 => x"81ff0bd4",
  1265 => x"0cd00870",
  1266 => x"8f2a7081",
  1267 => x"06515153",
  1268 => x"72f33872",
  1269 => x"d00c7580",
  1270 => x"d3a40c02",
  1271 => x"98050d04",
  1272 => x"02e8050d",
  1273 => x"77797b58",
  1274 => x"55558053",
  1275 => x"727625a3",
  1276 => x"38747081",
  1277 => x"055680f5",
  1278 => x"2d747081",
  1279 => x"055680f5",
  1280 => x"2d525271",
  1281 => x"712e8638",
  1282 => x"8151a895",
  1283 => x"04811353",
  1284 => x"a7ec0480",
  1285 => x"517080d3",
  1286 => x"a40c0298",
  1287 => x"050d0402",
  1288 => x"ec050d76",
  1289 => x"5574802e",
  1290 => x"80c2389a",
  1291 => x"1580e02d",
  1292 => x"51b6da2d",
  1293 => x"80d3a408",
  1294 => x"80d3a408",
  1295 => x"80dacc0c",
  1296 => x"80d3a408",
  1297 => x"545480da",
  1298 => x"a808802e",
  1299 => x"9a389415",
  1300 => x"80e02d51",
  1301 => x"b6da2d80",
  1302 => x"d3a40890",
  1303 => x"2b83fff0",
  1304 => x"0a067075",
  1305 => x"07515372",
  1306 => x"80dacc0c",
  1307 => x"80dacc08",
  1308 => x"5372802e",
  1309 => x"9d3880da",
  1310 => x"a008fe14",
  1311 => x"712980da",
  1312 => x"b4080580",
  1313 => x"dad00c70",
  1314 => x"842b80da",
  1315 => x"ac0c54a9",
  1316 => x"c00480da",
  1317 => x"b80880da",
  1318 => x"cc0c80da",
  1319 => x"bc0880da",
  1320 => x"d00c80da",
  1321 => x"a808802e",
  1322 => x"8b3880da",
  1323 => x"a008842b",
  1324 => x"53a9bb04",
  1325 => x"80dac008",
  1326 => x"842b5372",
  1327 => x"80daac0c",
  1328 => x"0294050d",
  1329 => x"0402d805",
  1330 => x"0d800b80",
  1331 => x"daa80c84",
  1332 => x"54a3ba2d",
  1333 => x"80d3a408",
  1334 => x"802e9738",
  1335 => x"80d49c52",
  1336 => x"8051a6bc",
  1337 => x"2d80d3a4",
  1338 => x"08802e86",
  1339 => x"38fe54a9",
  1340 => x"fa04ff14",
  1341 => x"54738024",
  1342 => x"d838738d",
  1343 => x"3880c9e4",
  1344 => x"5187f12d",
  1345 => x"7355afcf",
  1346 => x"04805681",
  1347 => x"0b80dad4",
  1348 => x"0c885380",
  1349 => x"c9f85280",
  1350 => x"d4d251a7",
  1351 => x"e02d80d3",
  1352 => x"a408762e",
  1353 => x"09810689",
  1354 => x"3880d3a4",
  1355 => x"0880dad4",
  1356 => x"0c885380",
  1357 => x"ca845280",
  1358 => x"d4ee51a7",
  1359 => x"e02d80d3",
  1360 => x"a4088938",
  1361 => x"80d3a408",
  1362 => x"80dad40c",
  1363 => x"80dad408",
  1364 => x"802e8181",
  1365 => x"3880d7e2",
  1366 => x"0b80f52d",
  1367 => x"80d7e30b",
  1368 => x"80f52d71",
  1369 => x"982b7190",
  1370 => x"2b0780d7",
  1371 => x"e40b80f5",
  1372 => x"2d70882b",
  1373 => x"720780d7",
  1374 => x"e50b80f5",
  1375 => x"2d710780",
  1376 => x"d89a0b80",
  1377 => x"f52d80d8",
  1378 => x"9b0b80f5",
  1379 => x"2d71882b",
  1380 => x"07535f54",
  1381 => x"525a5657",
  1382 => x"557381ab",
  1383 => x"aa2e0981",
  1384 => x"068e3875",
  1385 => x"51b6a92d",
  1386 => x"80d3a408",
  1387 => x"56abbe04",
  1388 => x"7382d4d5",
  1389 => x"2e883880",
  1390 => x"ca9051ac",
  1391 => x"8a0480d4",
  1392 => x"9c527551",
  1393 => x"a6bc2d80",
  1394 => x"d3a40855",
  1395 => x"80d3a408",
  1396 => x"802e83fb",
  1397 => x"38885380",
  1398 => x"ca845280",
  1399 => x"d4ee51a7",
  1400 => x"e02d80d3",
  1401 => x"a4088a38",
  1402 => x"810b80da",
  1403 => x"a80cac90",
  1404 => x"04885380",
  1405 => x"c9f85280",
  1406 => x"d4d251a7",
  1407 => x"e02d80d3",
  1408 => x"a408802e",
  1409 => x"8b3880ca",
  1410 => x"a45187f1",
  1411 => x"2dacef04",
  1412 => x"80d89a0b",
  1413 => x"80f52d54",
  1414 => x"7380d52e",
  1415 => x"09810680",
  1416 => x"ce3880d8",
  1417 => x"9b0b80f5",
  1418 => x"2d547381",
  1419 => x"aa2e0981",
  1420 => x"06bd3880",
  1421 => x"0b80d49c",
  1422 => x"0b80f52d",
  1423 => x"56547481",
  1424 => x"e92e8338",
  1425 => x"81547481",
  1426 => x"eb2e8c38",
  1427 => x"80557375",
  1428 => x"2e098106",
  1429 => x"82f93880",
  1430 => x"d4a70b80",
  1431 => x"f52d5574",
  1432 => x"8e3880d4",
  1433 => x"a80b80f5",
  1434 => x"2d547382",
  1435 => x"2e863880",
  1436 => x"55afcf04",
  1437 => x"80d4a90b",
  1438 => x"80f52d70",
  1439 => x"80daa00c",
  1440 => x"ff0580da",
  1441 => x"a40c80d4",
  1442 => x"aa0b80f5",
  1443 => x"2d80d4ab",
  1444 => x"0b80f52d",
  1445 => x"58760577",
  1446 => x"82802905",
  1447 => x"7080dab0",
  1448 => x"0c80d4ac",
  1449 => x"0b80f52d",
  1450 => x"7080dac4",
  1451 => x"0c80daa8",
  1452 => x"08595758",
  1453 => x"76802e81",
  1454 => x"b7388853",
  1455 => x"80ca8452",
  1456 => x"80d4ee51",
  1457 => x"a7e02d80",
  1458 => x"d3a40882",
  1459 => x"823880da",
  1460 => x"a0087084",
  1461 => x"2b80daac",
  1462 => x"0c7080da",
  1463 => x"c00c80d4",
  1464 => x"c10b80f5",
  1465 => x"2d80d4c0",
  1466 => x"0b80f52d",
  1467 => x"71828029",
  1468 => x"0580d4c2",
  1469 => x"0b80f52d",
  1470 => x"70848080",
  1471 => x"291280d4",
  1472 => x"c30b80f5",
  1473 => x"2d708180",
  1474 => x"0a291270",
  1475 => x"80dac80c",
  1476 => x"80dac408",
  1477 => x"712980da",
  1478 => x"b0080570",
  1479 => x"80dab40c",
  1480 => x"80d4c90b",
  1481 => x"80f52d80",
  1482 => x"d4c80b80",
  1483 => x"f52d7182",
  1484 => x"80290580",
  1485 => x"d4ca0b80",
  1486 => x"f52d7084",
  1487 => x"80802912",
  1488 => x"80d4cb0b",
  1489 => x"80f52d70",
  1490 => x"982b81f0",
  1491 => x"0a067205",
  1492 => x"7080dab8",
  1493 => x"0cfe117e",
  1494 => x"29770580",
  1495 => x"dabc0c52",
  1496 => x"59524354",
  1497 => x"5e515259",
  1498 => x"525d5759",
  1499 => x"57afc804",
  1500 => x"80d4ae0b",
  1501 => x"80f52d80",
  1502 => x"d4ad0b80",
  1503 => x"f52d7182",
  1504 => x"80290570",
  1505 => x"80daac0c",
  1506 => x"70a02983",
  1507 => x"ff057089",
  1508 => x"2a7080da",
  1509 => x"c00c80d4",
  1510 => x"b30b80f5",
  1511 => x"2d80d4b2",
  1512 => x"0b80f52d",
  1513 => x"71828029",
  1514 => x"057080da",
  1515 => x"c80c7b71",
  1516 => x"291e7080",
  1517 => x"dabc0c7d",
  1518 => x"80dab80c",
  1519 => x"730580da",
  1520 => x"b40c555e",
  1521 => x"51515555",
  1522 => x"8051a89f",
  1523 => x"2d815574",
  1524 => x"80d3a40c",
  1525 => x"02a8050d",
  1526 => x"0402ec05",
  1527 => x"0d767087",
  1528 => x"2c7180ff",
  1529 => x"06555654",
  1530 => x"80daa808",
  1531 => x"8a387388",
  1532 => x"2c7481ff",
  1533 => x"06545580",
  1534 => x"d49c5280",
  1535 => x"dab00815",
  1536 => x"51a6bc2d",
  1537 => x"80d3a408",
  1538 => x"5480d3a4",
  1539 => x"08802eb8",
  1540 => x"3880daa8",
  1541 => x"08802e9a",
  1542 => x"38728429",
  1543 => x"80d49c05",
  1544 => x"70085253",
  1545 => x"b6a92d80",
  1546 => x"d3a408f0",
  1547 => x"0a0653b0",
  1548 => x"c6047210",
  1549 => x"80d49c05",
  1550 => x"7080e02d",
  1551 => x"5253b6da",
  1552 => x"2d80d3a4",
  1553 => x"08537254",
  1554 => x"7380d3a4",
  1555 => x"0c029405",
  1556 => x"0d0402e0",
  1557 => x"050d7970",
  1558 => x"842c80da",
  1559 => x"d0080571",
  1560 => x"8f065255",
  1561 => x"53728a38",
  1562 => x"80d49c52",
  1563 => x"7351a6bc",
  1564 => x"2d72a029",
  1565 => x"80d49c05",
  1566 => x"54807480",
  1567 => x"f52d5653",
  1568 => x"74732e83",
  1569 => x"38815374",
  1570 => x"81e52e81",
  1571 => x"f4388170",
  1572 => x"74065458",
  1573 => x"72802e81",
  1574 => x"e8388b14",
  1575 => x"80f52d70",
  1576 => x"832a7906",
  1577 => x"5856769b",
  1578 => x"3880d1e8",
  1579 => x"08537289",
  1580 => x"387280d8",
  1581 => x"9c0b81b7",
  1582 => x"2d7680d1",
  1583 => x"e80c7353",
  1584 => x"b3830475",
  1585 => x"8f2e0981",
  1586 => x"0681b638",
  1587 => x"749f068d",
  1588 => x"2980d88f",
  1589 => x"11515381",
  1590 => x"1480f52d",
  1591 => x"73708105",
  1592 => x"5581b72d",
  1593 => x"831480f5",
  1594 => x"2d737081",
  1595 => x"055581b7",
  1596 => x"2d851480",
  1597 => x"f52d7370",
  1598 => x"81055581",
  1599 => x"b72d8714",
  1600 => x"80f52d73",
  1601 => x"70810555",
  1602 => x"81b72d89",
  1603 => x"1480f52d",
  1604 => x"73708105",
  1605 => x"5581b72d",
  1606 => x"8e1480f5",
  1607 => x"2d737081",
  1608 => x"055581b7",
  1609 => x"2d901480",
  1610 => x"f52d7370",
  1611 => x"81055581",
  1612 => x"b72d9214",
  1613 => x"80f52d73",
  1614 => x"70810555",
  1615 => x"81b72d94",
  1616 => x"1480f52d",
  1617 => x"73708105",
  1618 => x"5581b72d",
  1619 => x"961480f5",
  1620 => x"2d737081",
  1621 => x"055581b7",
  1622 => x"2d981480",
  1623 => x"f52d7370",
  1624 => x"81055581",
  1625 => x"b72d9c14",
  1626 => x"80f52d73",
  1627 => x"70810555",
  1628 => x"81b72d9e",
  1629 => x"1480f52d",
  1630 => x"7381b72d",
  1631 => x"7780d1e8",
  1632 => x"0c805372",
  1633 => x"80d3a40c",
  1634 => x"02a0050d",
  1635 => x"0402cc05",
  1636 => x"0d7e605e",
  1637 => x"5b800b80",
  1638 => x"dacc0880",
  1639 => x"dad00859",
  1640 => x"5d568059",
  1641 => x"80daac08",
  1642 => x"792e81de",
  1643 => x"38788f06",
  1644 => x"a0175754",
  1645 => x"73913880",
  1646 => x"d49c5276",
  1647 => x"51811757",
  1648 => x"a6bc2d80",
  1649 => x"d49c5680",
  1650 => x"7680f52d",
  1651 => x"56547474",
  1652 => x"2e833881",
  1653 => x"547481e5",
  1654 => x"2e81a338",
  1655 => x"81707506",
  1656 => x"555a7380",
  1657 => x"2e819738",
  1658 => x"8b1680f5",
  1659 => x"2d709806",
  1660 => x"59547780",
  1661 => x"e3388b53",
  1662 => x"7c527551",
  1663 => x"a7e02d80",
  1664 => x"d3a40880",
  1665 => x"f9389c16",
  1666 => x"0851b6a9",
  1667 => x"2d80d3a4",
  1668 => x"08841c0c",
  1669 => x"9a1680e0",
  1670 => x"2d51b6da",
  1671 => x"2d80d3a4",
  1672 => x"0880d3a4",
  1673 => x"08881d0c",
  1674 => x"80d3a408",
  1675 => x"555580da",
  1676 => x"a808802e",
  1677 => x"99389416",
  1678 => x"80e02d51",
  1679 => x"b6da2d80",
  1680 => x"d3a40890",
  1681 => x"2b83fff0",
  1682 => x"0a067016",
  1683 => x"51547388",
  1684 => x"1c0c777b",
  1685 => x"0cb4f904",
  1686 => x"73842a70",
  1687 => x"81065154",
  1688 => x"73802e9a",
  1689 => x"388b537c",
  1690 => x"527551a7",
  1691 => x"e02d80d3",
  1692 => x"a4088b38",
  1693 => x"7551a89f",
  1694 => x"2d7954b5",
  1695 => x"c6048119",
  1696 => x"5980daac",
  1697 => x"087926fe",
  1698 => x"a43880da",
  1699 => x"a808802e",
  1700 => x"b3387b51",
  1701 => x"afd92d80",
  1702 => x"d3a40880",
  1703 => x"d3a40880",
  1704 => x"fffffff8",
  1705 => x"06555c73",
  1706 => x"80ffffff",
  1707 => x"f82e9538",
  1708 => x"80d3a408",
  1709 => x"fe0580da",
  1710 => x"a0082980",
  1711 => x"dab40805",
  1712 => x"57b3a204",
  1713 => x"80547380",
  1714 => x"d3a40c02",
  1715 => x"b4050d04",
  1716 => x"02f4050d",
  1717 => x"74700881",
  1718 => x"05710c70",
  1719 => x"0880daa4",
  1720 => x"08065353",
  1721 => x"718f3888",
  1722 => x"130851af",
  1723 => x"d92d80d3",
  1724 => x"a4088814",
  1725 => x"0c810b80",
  1726 => x"d3a40c02",
  1727 => x"8c050d04",
  1728 => x"02f0050d",
  1729 => x"75881108",
  1730 => x"fe0580da",
  1731 => x"a0082980",
  1732 => x"dab40811",
  1733 => x"720880da",
  1734 => x"a4080605",
  1735 => x"79555354",
  1736 => x"54a6bc2d",
  1737 => x"0290050d",
  1738 => x"0402f405",
  1739 => x"0d747088",
  1740 => x"2a83fe80",
  1741 => x"06707298",
  1742 => x"2a077288",
  1743 => x"2b87fc80",
  1744 => x"80067398",
  1745 => x"2b81f00a",
  1746 => x"06717307",
  1747 => x"0780d3a4",
  1748 => x"0c565153",
  1749 => x"51028c05",
  1750 => x"0d0402f8",
  1751 => x"050d028e",
  1752 => x"0580f52d",
  1753 => x"74882b07",
  1754 => x"7083ffff",
  1755 => x"0680d3a4",
  1756 => x"0c510288",
  1757 => x"050d0402",
  1758 => x"ec050d76",
  1759 => x"787a5355",
  1760 => x"53815580",
  1761 => x"7125ae38",
  1762 => x"70527370",
  1763 => x"81055580",
  1764 => x"f52d7370",
  1765 => x"81055581",
  1766 => x"b72d7380",
  1767 => x"f52d5170",
  1768 => x"86387055",
  1769 => x"b7aa0474",
  1770 => x"8638a073",
  1771 => x"81b72dff",
  1772 => x"125271d6",
  1773 => x"38807381",
  1774 => x"b72d0294",
  1775 => x"050d0402",
  1776 => x"e8050d77",
  1777 => x"56807056",
  1778 => x"54737624",
  1779 => x"b63880da",
  1780 => x"ac08742e",
  1781 => x"ae387351",
  1782 => x"b0d22d80",
  1783 => x"d3a40880",
  1784 => x"d3a40809",
  1785 => x"81057080",
  1786 => x"d3a40807",
  1787 => x"9f2a7705",
  1788 => x"81175757",
  1789 => x"53537476",
  1790 => x"24893880",
  1791 => x"daac0874",
  1792 => x"26d43872",
  1793 => x"80d3a40c",
  1794 => x"0298050d",
  1795 => x"0402f005",
  1796 => x"0d80d3a0",
  1797 => x"081651b7",
  1798 => x"bf2d80d3",
  1799 => x"a408802e",
  1800 => x"9f388b53",
  1801 => x"80d3a408",
  1802 => x"5280d89c",
  1803 => x"51b6f72d",
  1804 => x"80dad808",
  1805 => x"5473802e",
  1806 => x"873880d8",
  1807 => x"9c51732d",
  1808 => x"0290050d",
  1809 => x"0402dc05",
  1810 => x"0d80705a",
  1811 => x"557480d3",
  1812 => x"a00825b4",
  1813 => x"3880daac",
  1814 => x"08752eac",
  1815 => x"387851b0",
  1816 => x"d22d80d3",
  1817 => x"a4080981",
  1818 => x"057080d3",
  1819 => x"a408079f",
  1820 => x"2a760581",
  1821 => x"1b5b5654",
  1822 => x"7480d3a0",
  1823 => x"08258938",
  1824 => x"80daac08",
  1825 => x"7926d638",
  1826 => x"80557880",
  1827 => x"daac0827",
  1828 => x"81db3878",
  1829 => x"51b0d22d",
  1830 => x"80d3a408",
  1831 => x"802e81ad",
  1832 => x"3880d3a4",
  1833 => x"088b0580",
  1834 => x"f52d7084",
  1835 => x"2a708106",
  1836 => x"77107884",
  1837 => x"2b80d89c",
  1838 => x"0b80f52d",
  1839 => x"5c5c5351",
  1840 => x"55567380",
  1841 => x"2e80cb38",
  1842 => x"7416822b",
  1843 => x"bb910b80",
  1844 => x"d1f4120c",
  1845 => x"54777531",
  1846 => x"1080dadc",
  1847 => x"11555690",
  1848 => x"74708105",
  1849 => x"5681b72d",
  1850 => x"a07481b7",
  1851 => x"2d7681ff",
  1852 => x"06811658",
  1853 => x"5473802e",
  1854 => x"8a389c53",
  1855 => x"80d89c52",
  1856 => x"ba8a048b",
  1857 => x"5380d3a4",
  1858 => x"085280da",
  1859 => x"de1651ba",
  1860 => x"c5047416",
  1861 => x"822bb88d",
  1862 => x"0b80d1f4",
  1863 => x"120c5476",
  1864 => x"81ff0681",
  1865 => x"16585473",
  1866 => x"802e8a38",
  1867 => x"9c5380d8",
  1868 => x"9c52babc",
  1869 => x"048b5380",
  1870 => x"d3a40852",
  1871 => x"77753110",
  1872 => x"80dadc05",
  1873 => x"517655b6",
  1874 => x"f72dbae2",
  1875 => x"04749029",
  1876 => x"75317010",
  1877 => x"80dadc05",
  1878 => x"515480d3",
  1879 => x"a4087481",
  1880 => x"b72d8119",
  1881 => x"59748b24",
  1882 => x"a338b98a",
  1883 => x"04749029",
  1884 => x"75317010",
  1885 => x"80dadc05",
  1886 => x"8c773157",
  1887 => x"51548074",
  1888 => x"81b72d9e",
  1889 => x"14ff1656",
  1890 => x"5474f338",
  1891 => x"02a4050d",
  1892 => x"0402fc05",
  1893 => x"0d80d3a0",
  1894 => x"081351b7",
  1895 => x"bf2d80d3",
  1896 => x"a408802e",
  1897 => x"893880d3",
  1898 => x"a40851a8",
  1899 => x"9f2d800b",
  1900 => x"80d3a00c",
  1901 => x"b8c52d93",
  1902 => x"8f2d0284",
  1903 => x"050d0402",
  1904 => x"f8050d73",
  1905 => x"5170fd2e",
  1906 => x"b13870fd",
  1907 => x"248a3870",
  1908 => x"fc2e80cd",
  1909 => x"38bcbb04",
  1910 => x"70fe2eb8",
  1911 => x"3870ff2e",
  1912 => x"09810680",
  1913 => x"d63880d3",
  1914 => x"a0085170",
  1915 => x"802e80cb",
  1916 => x"38ff1180",
  1917 => x"d3a00cbc",
  1918 => x"bb0480d3",
  1919 => x"a008f405",
  1920 => x"7080d3a0",
  1921 => x"0c517080",
  1922 => x"25b13880",
  1923 => x"0b80d3a0",
  1924 => x"0cbcbb04",
  1925 => x"80d3a008",
  1926 => x"810580d3",
  1927 => x"a00cbcbb",
  1928 => x"0480d3a0",
  1929 => x"088c1170",
  1930 => x"80d3a00c",
  1931 => x"525280da",
  1932 => x"ac087126",
  1933 => x"86387180",
  1934 => x"d3a00cb8",
  1935 => x"c52d938f",
  1936 => x"2d028805",
  1937 => x"0d0402fc",
  1938 => x"050d800b",
  1939 => x"80d3a00c",
  1940 => x"b8c52d91",
  1941 => x"fd2d80d3",
  1942 => x"a40880d3",
  1943 => x"900c80d1",
  1944 => x"ec5194b5",
  1945 => x"2d028405",
  1946 => x"0d0402f8",
  1947 => x"050d80d3",
  1948 => x"cc08bff9",
  1949 => x"ff068180",
  1950 => x"077080d3",
  1951 => x"cc0cfc0c",
  1952 => x"7351bcc6",
  1953 => x"2d028805",
  1954 => x"0d0402f8",
  1955 => x"050d80d3",
  1956 => x"cc08bffa",
  1957 => x"ff068280",
  1958 => x"077080d3",
  1959 => x"cc0cfc0c",
  1960 => x"7351bcc6",
  1961 => x"2d028805",
  1962 => x"0d0402f8",
  1963 => x"050d80d3",
  1964 => x"cc08bfff",
  1965 => x"ff068780",
  1966 => x"077080d3",
  1967 => x"cc0cfc0c",
  1968 => x"7351bcc6",
  1969 => x"2d028805",
  1970 => x"0d047180",
  1971 => x"dad80c04",
  1972 => x"00ffffff",
  1973 => x"ff00ffff",
  1974 => x"ffff00ff",
  1975 => x"ffffff00",
  1976 => x"436f6e74",
  1977 => x"696e7565",
  1978 => x"00000000",
  1979 => x"3d205a58",
  1980 => x"38312f5a",
  1981 => x"58383020",
  1982 => x"436f6e66",
  1983 => x"69677572",
  1984 => x"6174696f",
  1985 => x"6e203d00",
  1986 => x"3d3d3d3d",
  1987 => x"3d3d3d3d",
  1988 => x"3d3d3d3d",
  1989 => x"3d3d3d3d",
  1990 => x"3d3d3d3d",
  1991 => x"3d3d3d3d",
  1992 => x"3d3d3d00",
  1993 => x"4c6f7720",
  1994 => x"52414d3a",
  1995 => x"204f6666",
  1996 => x"2f384b42",
  1997 => x"00000000",
  1998 => x"51532043",
  1999 => x"4852533a",
  2000 => x"44697361",
  2001 => x"626c6564",
  2002 => x"2f456e61",
  2003 => x"626c6564",
  2004 => x"28463129",
  2005 => x"00000000",
  2006 => x"4348524f",
  2007 => x"4d413831",
  2008 => x"3a204469",
  2009 => x"7361626c",
  2010 => x"65642f45",
  2011 => x"6e61626c",
  2012 => x"65640000",
  2013 => x"496e7665",
  2014 => x"72736520",
  2015 => x"76696465",
  2016 => x"6f3a204f",
  2017 => x"66662f4f",
  2018 => x"6e000000",
  2019 => x"426c6163",
  2020 => x"6b20626f",
  2021 => x"72646572",
  2022 => x"3a204f66",
  2023 => x"662f4f6e",
  2024 => x"00000000",
  2025 => x"56696465",
  2026 => x"6f206672",
  2027 => x"65717565",
  2028 => x"6e63793a",
  2029 => x"20353048",
  2030 => x"7a2f3630",
  2031 => x"487a0000",
  2032 => x"476f2042",
  2033 => x"61636b00",
  2034 => x"536c6f77",
  2035 => x"206d6f64",
  2036 => x"65207370",
  2037 => x"6565643a",
  2038 => x"204f7269",
  2039 => x"67696e61",
  2040 => x"6c000000",
  2041 => x"536c6f77",
  2042 => x"206d6f64",
  2043 => x"65207370",
  2044 => x"6565643a",
  2045 => x"204e6f57",
  2046 => x"61697400",
  2047 => x"536c6f77",
  2048 => x"206d6f64",
  2049 => x"65207370",
  2050 => x"6565643a",
  2051 => x"20783200",
  2052 => x"536c6f77",
  2053 => x"206d6f64",
  2054 => x"65207370",
  2055 => x"6565643a",
  2056 => x"20783800",
  2057 => x"43485224",
  2058 => x"3132382f",
  2059 => x"5544473a",
  2060 => x"20313238",
  2061 => x"20436861",
  2062 => x"72730000",
  2063 => x"43485224",
  2064 => x"3132382f",
  2065 => x"5544473a",
  2066 => x"20363420",
  2067 => x"43686172",
  2068 => x"73000000",
  2069 => x"43485224",
  2070 => x"3132382f",
  2071 => x"5544473a",
  2072 => x"20446973",
  2073 => x"61626c65",
  2074 => x"64000000",
  2075 => x"4a6f7973",
  2076 => x"7469636b",
  2077 => x"3a204375",
  2078 => x"72736f72",
  2079 => x"00000000",
  2080 => x"4a6f7973",
  2081 => x"7469636b",
  2082 => x"3a205369",
  2083 => x"6e636c61",
  2084 => x"69720000",
  2085 => x"4a6f7973",
  2086 => x"7469636b",
  2087 => x"3a205a58",
  2088 => x"38310000",
  2089 => x"4d61696e",
  2090 => x"2052414d",
  2091 => x"3a203136",
  2092 => x"4b420000",
  2093 => x"4d61696e",
  2094 => x"2052414d",
  2095 => x"3a203332",
  2096 => x"4b420000",
  2097 => x"4d61696e",
  2098 => x"2052414d",
  2099 => x"3a203438",
  2100 => x"4b420000",
  2101 => x"4d61696e",
  2102 => x"2052414d",
  2103 => x"3a20314b",
  2104 => x"42000000",
  2105 => x"436f6d70",
  2106 => x"75746572",
  2107 => x"204d6f64",
  2108 => x"656c3a20",
  2109 => x"5a583831",
  2110 => x"00000000",
  2111 => x"436f6d70",
  2112 => x"75746572",
  2113 => x"204d6f64",
  2114 => x"656c3a20",
  2115 => x"5a583830",
  2116 => x"00000000",
  2117 => x"3d3d205a",
  2118 => x"5838312f",
  2119 => x"5a583830",
  2120 => x"20666f72",
  2121 => x"205a5844",
  2122 => x"4f53203d",
  2123 => x"3d000000",
  2124 => x"3d3d3d3d",
  2125 => x"3d3d3d3d",
  2126 => x"3d3d3d3d",
  2127 => x"3d3d3d3d",
  2128 => x"3d3d3d3d",
  2129 => x"3d3d3d3d",
  2130 => x"3d000000",
  2131 => x"52657365",
  2132 => x"74000000",
  2133 => x"4c6f6164",
  2134 => x"20546170",
  2135 => x"6520282e",
  2136 => x"70292010",
  2137 => x"00000000",
  2138 => x"4c6f6164",
  2139 => x"20546170",
  2140 => x"6520282e",
  2141 => x"6f292010",
  2142 => x"00000000",
  2143 => x"4c6f6164",
  2144 => x"20526f6d",
  2145 => x"2020282e",
  2146 => x"726f6d29",
  2147 => x"20100000",
  2148 => x"436f6e66",
  2149 => x"69677572",
  2150 => x"6174696f",
  2151 => x"6e206f70",
  2152 => x"74696f6e",
  2153 => x"73201000",
  2154 => x"4b657962",
  2155 => x"6f617264",
  2156 => x"2048656c",
  2157 => x"70000000",
  2158 => x"45786974",
  2159 => x"00000000",
  2160 => x"524f4d20",
  2161 => x"6c6f6164",
  2162 => x"696e6720",
  2163 => x"6661696c",
  2164 => x"65640000",
  2165 => x"4f4b0000",
  2166 => x"54617065",
  2167 => x"2066696c",
  2168 => x"65204c6f",
  2169 => x"61646564",
  2170 => x"2e000000",
  2171 => x"54797065",
  2172 => x"204c4f41",
  2173 => x"44202222",
  2174 => x"202b2045",
  2175 => x"4e544552",
  2176 => x"206f6e20",
  2177 => x"5a583831",
  2178 => x"00000000",
  2179 => x"5468656e",
  2180 => x"20707265",
  2181 => x"73732050",
  2182 => x"6c617920",
  2183 => x"616e6420",
  2184 => x"77616974",
  2185 => x"00000000",
  2186 => x"54686572",
  2187 => x"65206973",
  2188 => x"206e6f20",
  2189 => x"696d6167",
  2190 => x"65207768",
  2191 => x"656e206c",
  2192 => x"6f616469",
  2193 => x"6e670000",
  2194 => x"3d205a58",
  2195 => x"38312f5a",
  2196 => x"58383020",
  2197 => x"4b657962",
  2198 => x"6f617264",
  2199 => x"2048656c",
  2200 => x"70203d00",
  2201 => x"5363726f",
  2202 => x"6c6c204c",
  2203 => x"6f636b3a",
  2204 => x"20636861",
  2205 => x"6e676520",
  2206 => x"62657477",
  2207 => x"65656e00",
  2208 => x"52474220",
  2209 => x"616e6420",
  2210 => x"56474120",
  2211 => x"76696465",
  2212 => x"6f206d6f",
  2213 => x"64650000",
  2214 => x"4374726c",
  2215 => x"2b416c74",
  2216 => x"2b44656c",
  2217 => x"6574653a",
  2218 => x"20536f66",
  2219 => x"74205265",
  2220 => x"73657400",
  2221 => x"4374726c",
  2222 => x"2b416c74",
  2223 => x"2b426163",
  2224 => x"6b737061",
  2225 => x"63653a20",
  2226 => x"48617264",
  2227 => x"20726573",
  2228 => x"65740000",
  2229 => x"45736320",
  2230 => x"6f72206a",
  2231 => x"6f797374",
  2232 => x"69636b20",
  2233 => x"62742e32",
  2234 => x"3a20746f",
  2235 => x"2073686f",
  2236 => x"77000000",
  2237 => x"6f722068",
  2238 => x"69646520",
  2239 => x"74686520",
  2240 => x"6f707469",
  2241 => x"6f6e7320",
  2242 => x"6d656e75",
  2243 => x"2e000000",
  2244 => x"57415344",
  2245 => x"202f2063",
  2246 => x"7572736f",
  2247 => x"72206b65",
  2248 => x"7973202f",
  2249 => x"206a6f79",
  2250 => x"73746963",
  2251 => x"6b000000",
  2252 => x"746f2073",
  2253 => x"656c6563",
  2254 => x"74206d65",
  2255 => x"6e75206f",
  2256 => x"7074696f",
  2257 => x"6e2e0000",
  2258 => x"456e7465",
  2259 => x"72202f20",
  2260 => x"46697265",
  2261 => x"20746f20",
  2262 => x"63686f6f",
  2263 => x"7365206f",
  2264 => x"7074696f",
  2265 => x"6e2e0000",
  2266 => x"3d205a58",
  2267 => x"38312f5a",
  2268 => x"58383020",
  2269 => x"436f7265",
  2270 => x"20437265",
  2271 => x"64697473",
  2272 => x"20203d00",
  2273 => x"43686970",
  2274 => x"2d382063",
  2275 => x"6f726520",
  2276 => x"666f7220",
  2277 => x"5a58554e",
  2278 => x"4f2c2041",
  2279 => x"454f4e2c",
  2280 => x"00000000",
  2281 => x"5a58444f",
  2282 => x"5320616e",
  2283 => x"64205a58",
  2284 => x"444f532b",
  2285 => x"20626f61",
  2286 => x"7264732e",
  2287 => x"00000000",
  2288 => x"4f726967",
  2289 => x"696e616c",
  2290 => x"20636f72",
  2291 => x"65206279",
  2292 => x"3a000000",
  2293 => x"202d2043",
  2294 => x"61727374",
  2295 => x"656e2045",
  2296 => x"6c746f6e",
  2297 => x"20536f72",
  2298 => x"656e7365",
  2299 => x"6e200000",
  2300 => x"506f7274",
  2301 => x"206d6164",
  2302 => x"65206279",
  2303 => x"3a000000",
  2304 => x"202d2041",
  2305 => x"7a65736d",
  2306 => x"626f6700",
  2307 => x"202d2041",
  2308 => x"766c6978",
  2309 => x"41000000",
  2310 => x"496e6974",
  2311 => x"69616c69",
  2312 => x"7a696e67",
  2313 => x"20534420",
  2314 => x"63617264",
  2315 => x"0a000000",
  2316 => x"4c6f6164",
  2317 => x"696e6720",
  2318 => x"696e6974",
  2319 => x"69616c20",
  2320 => x"524f4d2e",
  2321 => x"2e2e0a00",
  2322 => x"5a583831",
  2323 => x"20202020",
  2324 => x"20202000",
  2325 => x"524f4d53",
  2326 => x"20202020",
  2327 => x"20202000",
  2328 => x"5a583858",
  2329 => x"20202020",
  2330 => x"524f4d00",
  2331 => x"4572726f",
  2332 => x"72204c6f",
  2333 => x"6164696e",
  2334 => x"6720524f",
  2335 => x"4d2e2e2e",
  2336 => x"0a000000",
  2337 => x"16200000",
  2338 => x"14200000",
  2339 => x"15200000",
  2340 => x"53442069",
  2341 => x"6e69742e",
  2342 => x"2e2e0a00",
  2343 => x"53442063",
  2344 => x"61726420",
  2345 => x"72657365",
  2346 => x"74206661",
  2347 => x"696c6564",
  2348 => x"210a0000",
  2349 => x"53444843",
  2350 => x"20657272",
  2351 => x"6f72210a",
  2352 => x"00000000",
  2353 => x"57726974",
  2354 => x"65206661",
  2355 => x"696c6564",
  2356 => x"0a000000",
  2357 => x"52656164",
  2358 => x"20666169",
  2359 => x"6c65640a",
  2360 => x"00000000",
  2361 => x"43617264",
  2362 => x"20696e69",
  2363 => x"74206661",
  2364 => x"696c6564",
  2365 => x"0a000000",
  2366 => x"46415431",
  2367 => x"36202020",
  2368 => x"00000000",
  2369 => x"46415433",
  2370 => x"32202020",
  2371 => x"00000000",
  2372 => x"4e6f2070",
  2373 => x"61727469",
  2374 => x"74696f6e",
  2375 => x"20736967",
  2376 => x"0a000000",
  2377 => x"42616420",
  2378 => x"70617274",
  2379 => x"0a000000",
  2380 => x"4261636b",
  2381 => x"00000000",
  2382 => x"00000002",
  2383 => x"00000002",
  2384 => x"00001eec",
  2385 => x"00000342",
  2386 => x"00000002",
  2387 => x"00001f08",
  2388 => x"00000342",
  2389 => x"00000003",
  2390 => x"00002628",
  2391 => x"00000002",
  2392 => x"00000003",
  2393 => x"00002618",
  2394 => x"00000004",
  2395 => x"00000001",
  2396 => x"00001f24",
  2397 => x"00000000",
  2398 => x"00000003",
  2399 => x"0000260c",
  2400 => x"00000003",
  2401 => x"00000001",
  2402 => x"00001f38",
  2403 => x"00000001",
  2404 => x"00000003",
  2405 => x"00002600",
  2406 => x"00000003",
  2407 => x"00000001",
  2408 => x"00001f58",
  2409 => x"00000002",
  2410 => x"00000001",
  2411 => x"00001f74",
  2412 => x"00000003",
  2413 => x"00000001",
  2414 => x"00001f8c",
  2415 => x"00000004",
  2416 => x"00000003",
  2417 => x"000025f0",
  2418 => x"00000003",
  2419 => x"00000001",
  2420 => x"00001fa4",
  2421 => x"00000005",
  2422 => x"00000004",
  2423 => x"00001fc0",
  2424 => x"000029d0",
  2425 => x"00000000",
  2426 => x"00000000",
  2427 => x"00000000",
  2428 => x"00001fc8",
  2429 => x"00001fe4",
  2430 => x"00001ffc",
  2431 => x"00002010",
  2432 => x"00002024",
  2433 => x"0000203c",
  2434 => x"00002054",
  2435 => x"0000206c",
  2436 => x"00002080",
  2437 => x"00002094",
  2438 => x"000020a4",
  2439 => x"000020b4",
  2440 => x"000020c4",
  2441 => x"000020d4",
  2442 => x"000020e4",
  2443 => x"000020fc",
  2444 => x"00000002",
  2445 => x"00002114",
  2446 => x"00000343",
  2447 => x"00000002",
  2448 => x"00002130",
  2449 => x"00000343",
  2450 => x"00000002",
  2451 => x"0000214c",
  2452 => x"00000386",
  2453 => x"00000002",
  2454 => x"00002154",
  2455 => x"00001e6a",
  2456 => x"00000002",
  2457 => x"00002168",
  2458 => x"00001e8a",
  2459 => x"00000002",
  2460 => x"0000217c",
  2461 => x"00001eaa",
  2462 => x"00000002",
  2463 => x"00002190",
  2464 => x"00000353",
  2465 => x"00000002",
  2466 => x"000021a8",
  2467 => x"00000363",
  2468 => x"00000002",
  2469 => x"000021b8",
  2470 => x"0000091a",
  2471 => x"00000000",
  2472 => x"00000000",
  2473 => x"00000000",
  2474 => x"00000004",
  2475 => x"000021c0",
  2476 => x"000026a8",
  2477 => x"00000004",
  2478 => x"000021d4",
  2479 => x"000029d0",
  2480 => x"00000000",
  2481 => x"00000000",
  2482 => x"00000000",
  2483 => x"00000004",
  2484 => x"000021d8",
  2485 => x"000026cc",
  2486 => x"00000004",
  2487 => x"000021ec",
  2488 => x"000026cc",
  2489 => x"00000004",
  2490 => x"0000220c",
  2491 => x"000026cc",
  2492 => x"00000004",
  2493 => x"00002228",
  2494 => x"000026cc",
  2495 => x"00000004",
  2496 => x"000024c0",
  2497 => x"000026cc",
  2498 => x"00000004",
  2499 => x"00001ee0",
  2500 => x"000029d0",
  2501 => x"00000000",
  2502 => x"00000000",
  2503 => x"00000000",
  2504 => x"00000002",
  2505 => x"00002248",
  2506 => x"00000342",
  2507 => x"00000002",
  2508 => x"00001f08",
  2509 => x"00000342",
  2510 => x"00000002",
  2511 => x"00002264",
  2512 => x"00000342",
  2513 => x"00000002",
  2514 => x"00002280",
  2515 => x"00000342",
  2516 => x"00000002",
  2517 => x"00002298",
  2518 => x"00000342",
  2519 => x"00000002",
  2520 => x"000022b4",
  2521 => x"00000342",
  2522 => x"00000002",
  2523 => x"000022d4",
  2524 => x"00000342",
  2525 => x"00000002",
  2526 => x"000022f4",
  2527 => x"00000342",
  2528 => x"00000002",
  2529 => x"00002310",
  2530 => x"00000342",
  2531 => x"00000002",
  2532 => x"00002330",
  2533 => x"00000342",
  2534 => x"00000002",
  2535 => x"00002348",
  2536 => x"00000342",
  2537 => x"00000002",
  2538 => x"000024c0",
  2539 => x"00000342",
  2540 => x"00000004",
  2541 => x"000021d4",
  2542 => x"000029d0",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000002",
  2547 => x"00002368",
  2548 => x"00000342",
  2549 => x"00000002",
  2550 => x"00001f08",
  2551 => x"00000342",
  2552 => x"00000002",
  2553 => x"00002384",
  2554 => x"00000342",
  2555 => x"00000002",
  2556 => x"000023a4",
  2557 => x"00000342",
  2558 => x"00000002",
  2559 => x"000024c0",
  2560 => x"00000342",
  2561 => x"00000002",
  2562 => x"000023c0",
  2563 => x"00000342",
  2564 => x"00000002",
  2565 => x"000023d4",
  2566 => x"00000342",
  2567 => x"00000002",
  2568 => x"000024c0",
  2569 => x"00000342",
  2570 => x"00000002",
  2571 => x"000023f0",
  2572 => x"00000342",
  2573 => x"00000002",
  2574 => x"00002400",
  2575 => x"00000342",
  2576 => x"00000002",
  2577 => x"0000240c",
  2578 => x"00000342",
  2579 => x"00000002",
  2580 => x"000024c0",
  2581 => x"00000342",
  2582 => x"00000004",
  2583 => x"000021d4",
  2584 => x"000029d0",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000006",
  2607 => x"00000043",
  2608 => x"00000042",
  2609 => x"0000003b",
  2610 => x"0000004b",
  2611 => x"0000007e",
  2612 => x"00000003",
  2613 => x"0000000b",
  2614 => x"00000083",
  2615 => x"00000023",
  2616 => x"0000007e",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000002",
  2620 => x"00002d5c",
  2621 => x"00001c0d",
  2622 => x"00000002",
  2623 => x"00002d7a",
  2624 => x"00001c0d",
  2625 => x"00000002",
  2626 => x"00002d98",
  2627 => x"00001c0d",
  2628 => x"00000002",
  2629 => x"00002db6",
  2630 => x"00001c0d",
  2631 => x"00000002",
  2632 => x"00002dd4",
  2633 => x"00001c0d",
  2634 => x"00000002",
  2635 => x"00002df2",
  2636 => x"00001c0d",
  2637 => x"00000002",
  2638 => x"00002e10",
  2639 => x"00001c0d",
  2640 => x"00000002",
  2641 => x"00002e2e",
  2642 => x"00001c0d",
  2643 => x"00000002",
  2644 => x"00002e4c",
  2645 => x"00001c0d",
  2646 => x"00000002",
  2647 => x"00002e6a",
  2648 => x"00001c0d",
  2649 => x"00000002",
  2650 => x"00002e88",
  2651 => x"00001c0d",
  2652 => x"00000002",
  2653 => x"00002ea6",
  2654 => x"00001c0d",
  2655 => x"00000002",
  2656 => x"00002ec4",
  2657 => x"00001c0d",
  2658 => x"00000004",
  2659 => x"00002530",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00001dbf",
  2664 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

