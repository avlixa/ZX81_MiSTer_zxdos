-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d5",
     9 => x"d4080b0b",
    10 => x"80d5d808",
    11 => x"0b0b80d5",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d5dc0c0b",
    16 => x"0b80d5d8",
    17 => x"0c0b0b80",
    18 => x"d5d40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbef0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d5d470",
    57 => x"80e09427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518add",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d5",
    65 => x"e40c9f0b",
    66 => x"80d5e80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d5e808ff",
    70 => x"0580d5e8",
    71 => x"0c80d5e8",
    72 => x"088025e8",
    73 => x"3880d5e4",
    74 => x"08ff0580",
    75 => x"d5e40c80",
    76 => x"d5e40880",
    77 => x"25d03880",
    78 => x"0b80d5e8",
    79 => x"0c800b80",
    80 => x"d5e40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d5e408",
   100 => x"25913882",
   101 => x"c82d80d5",
   102 => x"e408ff05",
   103 => x"80d5e40c",
   104 => x"838a0480",
   105 => x"d5e40880",
   106 => x"d5e80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d5e408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d5e80881",
   116 => x"0580d5e8",
   117 => x"0c80d5e8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d5e8",
   121 => x"0c80d5e4",
   122 => x"08810580",
   123 => x"d5e40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d5",
   128 => x"e8088105",
   129 => x"80d5e80c",
   130 => x"80d5e808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d5e8",
   134 => x"0c80d5e4",
   135 => x"08810580",
   136 => x"d5e40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d5ec0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d5ec0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d5",
   177 => x"ec088407",
   178 => x"80d5ec0c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5483f474",
   182 => x"258f3883",
   183 => x"0b0b0b80",
   184 => x"cbec0c82",
   185 => x"985385f3",
   186 => x"04810b0b",
   187 => x"0b80cbec",
   188 => x"0ca8530b",
   189 => x"0b80cbec",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0c747431",
   193 => x"ffb005ff",
   194 => x"1271712c",
   195 => x"ff941970",
   196 => x"9f2a1170",
   197 => x"812c80d5",
   198 => x"ec085255",
   199 => x"51525652",
   200 => x"53517680",
   201 => x"2e853870",
   202 => x"81075170",
   203 => x"f6940c72",
   204 => x"098105f6",
   205 => x"800c7109",
   206 => x"8105f684",
   207 => x"0c029405",
   208 => x"0d040402",
   209 => x"fc050d80",
   210 => x"d1f85195",
   211 => x"c52d0284",
   212 => x"050d0402",
   213 => x"fc050d80",
   214 => x"cbf05195",
   215 => x"c52d0284",
   216 => x"050d0402",
   217 => x"fc050d80",
   218 => x"d0d05195",
   219 => x"c52d0284",
   220 => x"050d0402",
   221 => x"fc050d81",
   222 => x"808051c0",
   223 => x"115170fb",
   224 => x"38028405",
   225 => x"0d047181",
   226 => x"2e098106",
   227 => x"893881c3",
   228 => x"0bec0c87",
   229 => x"9a04830b",
   230 => x"ec0c86f3",
   231 => x"2d820bec",
   232 => x"0c049388",
   233 => x"2d80d5d4",
   234 => x"0880d0c0",
   235 => x"0c93882d",
   236 => x"80d5d408",
   237 => x"80cfec0c",
   238 => x"93882d80",
   239 => x"d5d40880",
   240 => x"d3900c93",
   241 => x"882d80d5",
   242 => x"d40880d1",
   243 => x"e80c9388",
   244 => x"2d80d5d4",
   245 => x"0880cd94",
   246 => x"0c0402fc",
   247 => x"050d84bf",
   248 => x"5186f32d",
   249 => x"ff115170",
   250 => x"8025f638",
   251 => x"0284050d",
   252 => x"0402f405",
   253 => x"0d745372",
   254 => x"70810554",
   255 => x"80f52d52",
   256 => x"71802e89",
   257 => x"38715183",
   258 => x"842d87f7",
   259 => x"04810b80",
   260 => x"d5d40c02",
   261 => x"8c050d04",
   262 => x"02dc050d",
   263 => x"800b80cd",
   264 => x"e4085459",
   265 => x"72822e89",
   266 => x"3872832e",
   267 => x"963888d5",
   268 => x"0480d5fc",
   269 => x"08bffaff",
   270 => x"06828007",
   271 => x"80d5fc0c",
   272 => x"88e40480",
   273 => x"d5fc08bf",
   274 => x"ffff0687",
   275 => x"800780d5",
   276 => x"fc0c88e4",
   277 => x"0480d5fc",
   278 => x"08bff9ff",
   279 => x"06818007",
   280 => x"80d5fc0c",
   281 => x"80d5fc08",
   282 => x"fc0c8184",
   283 => x"0bec0c7a",
   284 => x"5280d5f0",
   285 => x"51b49b2d",
   286 => x"80d5d408",
   287 => x"802e819d",
   288 => x"3880d5f4",
   289 => x"08548056",
   290 => x"73852e09",
   291 => x"81068a38",
   292 => x"840bec0c",
   293 => x"81538aa5",
   294 => x"0473f80c",
   295 => x"81a40bec",
   296 => x"0c87da2d",
   297 => x"75ff1557",
   298 => x"5875802e",
   299 => x"8b388118",
   300 => x"76812a57",
   301 => x"5889a904",
   302 => x"f7185881",
   303 => x"59807425",
   304 => x"80d738a4",
   305 => x"0bec0c77",
   306 => x"52755184",
   307 => x"a82d80d6",
   308 => x"cc5280d5",
   309 => x"f051b78e",
   310 => x"2d80d5d4",
   311 => x"08802ea0",
   312 => x"3880d6cc",
   313 => x"5783fc55",
   314 => x"76708405",
   315 => x"5808e80c",
   316 => x"fc155574",
   317 => x"8025f138",
   318 => x"81a40bec",
   319 => x"0c8a8804",
   320 => x"80d5d408",
   321 => x"59848054",
   322 => x"80d5f051",
   323 => x"b6de2dfc",
   324 => x"80148117",
   325 => x"575489bd",
   326 => x"04840bec",
   327 => x"0c80d5f4",
   328 => x"08f80c78",
   329 => x"537280d5",
   330 => x"d40c02a4",
   331 => x"050d0402",
   332 => x"f8050d73",
   333 => x"5188982d",
   334 => x"80d5d408",
   335 => x"5280d5d4",
   336 => x"08802e88",
   337 => x"3880cffc",
   338 => x"518ad004",
   339 => x"80cfd851",
   340 => x"95c52d71",
   341 => x"80d5d40c",
   342 => x"0288050d",
   343 => x"0402f005",
   344 => x"0d800b80",
   345 => x"d5fc0c81",
   346 => x"5187862d",
   347 => x"80518786",
   348 => x"2d840bec",
   349 => x"0c92d82d",
   350 => x"8f832d81",
   351 => x"f92d8352",
   352 => x"92bb2d81",
   353 => x"51858d2d",
   354 => x"ff125271",
   355 => x"8025f138",
   356 => x"80c40bec",
   357 => x"0c80c9c0",
   358 => x"5187f12d",
   359 => x"aad32d80",
   360 => x"d5d40880",
   361 => x"2e83c538",
   362 => x"81840bec",
   363 => x"0c80c9d8",
   364 => x"5187f12d",
   365 => x"80d5fc08",
   366 => x"bfffff06",
   367 => x"87800770",
   368 => x"80d5fc0c",
   369 => x"fc0c80c9",
   370 => x"f0518898",
   371 => x"2d80d5d4",
   372 => x"08802e80",
   373 => x"cc3880c9",
   374 => x"fc518898",
   375 => x"2d80d5d4",
   376 => x"08802ebd",
   377 => x"3880ca88",
   378 => x"5188982d",
   379 => x"80d5d408",
   380 => x"5280d5d4",
   381 => x"08973880",
   382 => x"ca945187",
   383 => x"f12d80ca",
   384 => x"ac518898",
   385 => x"2d715187",
   386 => x"862d8ca8",
   387 => x"0480caac",
   388 => x"5188982d",
   389 => x"80518786",
   390 => x"2d805185",
   391 => x"8d2d8ca8",
   392 => x"0480ca94",
   393 => x"5187f12d",
   394 => x"840bec0c",
   395 => x"8aaf51be",
   396 => x"ea2d80d5",
   397 => x"fc0880d3",
   398 => x"e80c80d5",
   399 => x"fc08fc0c",
   400 => x"80d6ac08",
   401 => x"882a7081",
   402 => x"06515271",
   403 => x"802e8c38",
   404 => x"80cee00b",
   405 => x"80d6800c",
   406 => x"8ce30480",
   407 => x"cde80b80",
   408 => x"d6800c80",
   409 => x"d6800851",
   410 => x"95c52d80",
   411 => x"5187a22d",
   412 => x"830b80d6",
   413 => x"c00c9391",
   414 => x"2d805185",
   415 => x"8d2d93a5",
   416 => x"2d8f8f2d",
   417 => x"95d82d80",
   418 => x"cc900b80",
   419 => x"f52d80cc",
   420 => x"9c0b80f5",
   421 => x"2d718a2b",
   422 => x"718b2b07",
   423 => x"80ccb40b",
   424 => x"80f52d70",
   425 => x"8d2b7207",
   426 => x"80cccc0b",
   427 => x"80f52d70",
   428 => x"8e2b7207",
   429 => x"80ccfc0b",
   430 => x"80f52d70",
   431 => x"912b7207",
   432 => x"7080d5fc",
   433 => x"0c80d3e8",
   434 => x"08708106",
   435 => x"54525354",
   436 => x"52545253",
   437 => x"54555371",
   438 => x"802e8838",
   439 => x"73810780",
   440 => x"d5fc0c72",
   441 => x"812a7081",
   442 => x"06515271",
   443 => x"802e8b38",
   444 => x"80d5fc08",
   445 => x"820780d5",
   446 => x"fc0c7282",
   447 => x"2a708106",
   448 => x"51527180",
   449 => x"2e8b3880",
   450 => x"d5fc0884",
   451 => x"0780d5fc",
   452 => x"0c72832a",
   453 => x"70810651",
   454 => x"5271802e",
   455 => x"8b3880d5",
   456 => x"fc088807",
   457 => x"80d5fc0c",
   458 => x"72842a70",
   459 => x"81065152",
   460 => x"71802e8b",
   461 => x"3880d5fc",
   462 => x"08900780",
   463 => x"d5fc0c72",
   464 => x"852a7081",
   465 => x"06515271",
   466 => x"802e8b38",
   467 => x"80d5fc08",
   468 => x"a00780d5",
   469 => x"fc0c80d5",
   470 => x"fc08fc0c",
   471 => x"865280d5",
   472 => x"d4088338",
   473 => x"845271ec",
   474 => x"0c8d8104",
   475 => x"800b80d5",
   476 => x"d40c0290",
   477 => x"050d0471",
   478 => x"980c04ff",
   479 => x"b00880d5",
   480 => x"d40c0481",
   481 => x"0bffb00c",
   482 => x"04800bff",
   483 => x"b00c0402",
   484 => x"f4050d90",
   485 => x"9d0480d5",
   486 => x"d40881f0",
   487 => x"2e098106",
   488 => x"8a38810b",
   489 => x"80d3e00c",
   490 => x"909d0480",
   491 => x"d5d40881",
   492 => x"e02e0981",
   493 => x"068a3881",
   494 => x"0b80d3e4",
   495 => x"0c909d04",
   496 => x"80d5d408",
   497 => x"5280d3e4",
   498 => x"08802e89",
   499 => x"3880d5d4",
   500 => x"08818005",
   501 => x"5271842c",
   502 => x"728f0653",
   503 => x"5380d3e0",
   504 => x"08802e9a",
   505 => x"38728429",
   506 => x"80d3a005",
   507 => x"72138171",
   508 => x"2b700973",
   509 => x"0806730c",
   510 => x"51535390",
   511 => x"91047284",
   512 => x"2980d3a0",
   513 => x"05721383",
   514 => x"712b7208",
   515 => x"07720c53",
   516 => x"53800b80",
   517 => x"d3e40c80",
   518 => x"0b80d3e0",
   519 => x"0c80d684",
   520 => x"5191a42d",
   521 => x"80d5d408",
   522 => x"ff24feea",
   523 => x"38800b80",
   524 => x"d5d40c02",
   525 => x"8c050d04",
   526 => x"02f8050d",
   527 => x"80d3a052",
   528 => x"8f518072",
   529 => x"70840554",
   530 => x"0cff1151",
   531 => x"708025f2",
   532 => x"38028805",
   533 => x"0d0402f0",
   534 => x"050d7551",
   535 => x"8f892d70",
   536 => x"822cfc06",
   537 => x"80d3a011",
   538 => x"72109e06",
   539 => x"71087072",
   540 => x"2a708306",
   541 => x"82742b70",
   542 => x"09740676",
   543 => x"0c545156",
   544 => x"57535153",
   545 => x"8f832d71",
   546 => x"80d5d40c",
   547 => x"0290050d",
   548 => x"0402fc05",
   549 => x"0d725180",
   550 => x"710c800b",
   551 => x"84120c02",
   552 => x"84050d04",
   553 => x"02f0050d",
   554 => x"75700884",
   555 => x"12085353",
   556 => x"53ff5471",
   557 => x"712ea838",
   558 => x"8f892d84",
   559 => x"13087084",
   560 => x"29148811",
   561 => x"70087081",
   562 => x"ff068418",
   563 => x"08811187",
   564 => x"06841a0c",
   565 => x"53515551",
   566 => x"51518f83",
   567 => x"2d715473",
   568 => x"80d5d40c",
   569 => x"0290050d",
   570 => x"0402f405",
   571 => x"0d8f892d",
   572 => x"e008708b",
   573 => x"2a708106",
   574 => x"51525370",
   575 => x"802ea138",
   576 => x"80d68408",
   577 => x"70842980",
   578 => x"d68c0574",
   579 => x"81ff0671",
   580 => x"0c515180",
   581 => x"d6840881",
   582 => x"11870680",
   583 => x"d6840c51",
   584 => x"728c2c83",
   585 => x"ff0680d6",
   586 => x"ac0c800b",
   587 => x"80d6b00c",
   588 => x"8efb2d8f",
   589 => x"832d028c",
   590 => x"050d0402",
   591 => x"fc050d8f",
   592 => x"892d810b",
   593 => x"80d6b00c",
   594 => x"8f832d80",
   595 => x"d6b00851",
   596 => x"70f93802",
   597 => x"84050d04",
   598 => x"02fc050d",
   599 => x"80d68451",
   600 => x"91912d90",
   601 => x"b82d91e9",
   602 => x"518ef72d",
   603 => x"0284050d",
   604 => x"0402fc05",
   605 => x"0d8fcf51",
   606 => x"86f32dff",
   607 => x"11517080",
   608 => x"25f63802",
   609 => x"84050d04",
   610 => x"80d6b808",
   611 => x"80d5d40c",
   612 => x"0402fc05",
   613 => x"0d810b80",
   614 => x"d4940c81",
   615 => x"51858d2d",
   616 => x"0284050d",
   617 => x"0402f805",
   618 => x"0d93af04",
   619 => x"8f8f2d80",
   620 => x"da5190d6",
   621 => x"2d80d5d4",
   622 => x"08810652",
   623 => x"71ee3880",
   624 => x"d4900851",
   625 => x"90d62d80",
   626 => x"d5d40881",
   627 => x"065271dc",
   628 => x"38835190",
   629 => x"d62d80d5",
   630 => x"d4088106",
   631 => x"5271cd38",
   632 => x"7180d494",
   633 => x"0c715185",
   634 => x"8d2d0288",
   635 => x"050d0402",
   636 => x"ec050d76",
   637 => x"54805287",
   638 => x"0b881580",
   639 => x"f52d5653",
   640 => x"74722483",
   641 => x"38a05372",
   642 => x"5183842d",
   643 => x"81128b15",
   644 => x"80f52d54",
   645 => x"52727225",
   646 => x"de380294",
   647 => x"050d0402",
   648 => x"f0050d80",
   649 => x"d6b80854",
   650 => x"81f92d80",
   651 => x"0b80d6bc",
   652 => x"0c730880",
   653 => x"2e818938",
   654 => x"820b80d5",
   655 => x"e80c80d6",
   656 => x"bc088f06",
   657 => x"80d5e40c",
   658 => x"73085271",
   659 => x"832e9638",
   660 => x"71832689",
   661 => x"3871812e",
   662 => x"b03895a9",
   663 => x"0471852e",
   664 => x"a03895a9",
   665 => x"04881480",
   666 => x"f52d8415",
   667 => x"0880cab8",
   668 => x"53545287",
   669 => x"f12d7184",
   670 => x"29137008",
   671 => x"525295ad",
   672 => x"04735193",
   673 => x"ef2d95a9",
   674 => x"0480d3e8",
   675 => x"08881508",
   676 => x"2c708106",
   677 => x"51527180",
   678 => x"2e883880",
   679 => x"cabc5195",
   680 => x"a60480ca",
   681 => x"c05187f1",
   682 => x"2d841408",
   683 => x"5187f12d",
   684 => x"80d6bc08",
   685 => x"810580d6",
   686 => x"bc0c8c14",
   687 => x"5494b104",
   688 => x"0290050d",
   689 => x"047180d6",
   690 => x"b80c949f",
   691 => x"2d80d6bc",
   692 => x"08ff0580",
   693 => x"d6c00c04",
   694 => x"02e8050d",
   695 => x"80d6b808",
   696 => x"80d6c408",
   697 => x"57558351",
   698 => x"90d62d80",
   699 => x"d5d40883",
   700 => x"06527180",
   701 => x"2ea53895",
   702 => x"fd048f8f",
   703 => x"2d835190",
   704 => x"d62d80d5",
   705 => x"d4088106",
   706 => x"5271ef38",
   707 => x"80d49408",
   708 => x"81327080",
   709 => x"d4940c51",
   710 => x"858d2d80",
   711 => x"0b80d6b4",
   712 => x"0c8c5190",
   713 => x"d62d80d5",
   714 => x"d408812a",
   715 => x"70810651",
   716 => x"5271802e",
   717 => x"80d13880",
   718 => x"d3ec0880",
   719 => x"d4800880",
   720 => x"d3ec0c80",
   721 => x"d4800c80",
   722 => x"d3f00880",
   723 => x"d4840880",
   724 => x"d3f00c80",
   725 => x"d4840c80",
   726 => x"d3f40880",
   727 => x"d4880880",
   728 => x"d3f40c80",
   729 => x"d4880c80",
   730 => x"d3f80880",
   731 => x"d48c0880",
   732 => x"d3f80c80",
   733 => x"d48c0c80",
   734 => x"d3fc0880",
   735 => x"d4900880",
   736 => x"d3fc0c80",
   737 => x"d4900c80",
   738 => x"d6ac08a0",
   739 => x"06528072",
   740 => x"25963892",
   741 => x"f12d8f8f",
   742 => x"2d80d494",
   743 => x"08813270",
   744 => x"80d4940c",
   745 => x"51858d2d",
   746 => x"80d49408",
   747 => x"82ef3880",
   748 => x"d4800851",
   749 => x"90d62d80",
   750 => x"d5d40880",
   751 => x"2e8b3880",
   752 => x"d6b40881",
   753 => x"0780d6b4",
   754 => x"0c80d484",
   755 => x"085190d6",
   756 => x"2d80d5d4",
   757 => x"08802e8b",
   758 => x"3880d6b4",
   759 => x"08820780",
   760 => x"d6b40c80",
   761 => x"d4880851",
   762 => x"90d62d80",
   763 => x"d5d40880",
   764 => x"2e8b3880",
   765 => x"d6b40884",
   766 => x"0780d6b4",
   767 => x"0c80d48c",
   768 => x"085190d6",
   769 => x"2d80d5d4",
   770 => x"08802e8b",
   771 => x"3880d6b4",
   772 => x"08880780",
   773 => x"d6b40c80",
   774 => x"d4900851",
   775 => x"90d62d80",
   776 => x"d5d40880",
   777 => x"2e8b3880",
   778 => x"d6b40890",
   779 => x"0780d6b4",
   780 => x"0c80d3ec",
   781 => x"085190d6",
   782 => x"2d80d5d4",
   783 => x"08802e8c",
   784 => x"3880d6b4",
   785 => x"08828007",
   786 => x"80d6b40c",
   787 => x"80d3f008",
   788 => x"5190d62d",
   789 => x"80d5d408",
   790 => x"802e8c38",
   791 => x"80d6b408",
   792 => x"84800780",
   793 => x"d6b40c80",
   794 => x"d3f40851",
   795 => x"90d62d80",
   796 => x"d5d40880",
   797 => x"2e8c3880",
   798 => x"d6b40888",
   799 => x"800780d6",
   800 => x"b40c80d3",
   801 => x"f8085190",
   802 => x"d62d80d5",
   803 => x"d408802e",
   804 => x"8c3880d6",
   805 => x"b4089080",
   806 => x"0780d6b4",
   807 => x"0c80d3fc",
   808 => x"085190d6",
   809 => x"2d80d5d4",
   810 => x"08802e8c",
   811 => x"3880d6b4",
   812 => x"08a08007",
   813 => x"80d6b40c",
   814 => x"945190d6",
   815 => x"2d80d5d4",
   816 => x"08529151",
   817 => x"90d62d71",
   818 => x"80d5d408",
   819 => x"065280e6",
   820 => x"5190d62d",
   821 => x"7180d5d4",
   822 => x"08065271",
   823 => x"802e8d38",
   824 => x"80d6b408",
   825 => x"84808007",
   826 => x"80d6b40c",
   827 => x"80fe5190",
   828 => x"d62d80d5",
   829 => x"d4085287",
   830 => x"5190d62d",
   831 => x"7180d5d4",
   832 => x"08075271",
   833 => x"802e8d38",
   834 => x"80d6b408",
   835 => x"88808007",
   836 => x"80d6b40c",
   837 => x"80d6b408",
   838 => x"ed0ca2a8",
   839 => x"04945190",
   840 => x"d62d80d5",
   841 => x"d4085291",
   842 => x"5190d62d",
   843 => x"7180d5d4",
   844 => x"08065280",
   845 => x"e65190d6",
   846 => x"2d7180d5",
   847 => x"d4080652",
   848 => x"71802e8d",
   849 => x"3880d6b4",
   850 => x"08848080",
   851 => x"0780d6b4",
   852 => x"0c80fe51",
   853 => x"90d62d80",
   854 => x"d5d40852",
   855 => x"875190d6",
   856 => x"2d7180d5",
   857 => x"d4080752",
   858 => x"71802e8d",
   859 => x"3880d6b4",
   860 => x"08888080",
   861 => x"0780d6b4",
   862 => x"0c80d6b4",
   863 => x"08ed0c81",
   864 => x"f55190d6",
   865 => x"2d80d5d4",
   866 => x"08812a70",
   867 => x"81065152",
   868 => x"71a43880",
   869 => x"d4800851",
   870 => x"90d62d80",
   871 => x"d5d40881",
   872 => x"2a708106",
   873 => x"5152718e",
   874 => x"3880d6ac",
   875 => x"08810652",
   876 => x"80722580",
   877 => x"c23880d6",
   878 => x"ac088106",
   879 => x"52807225",
   880 => x"843892f1",
   881 => x"2d80d6c0",
   882 => x"08527180",
   883 => x"2e8a38ff",
   884 => x"1280d6c0",
   885 => x"0c9bf704",
   886 => x"80d6bc08",
   887 => x"1080d6bc",
   888 => x"08057084",
   889 => x"29165152",
   890 => x"88120880",
   891 => x"2e8938ff",
   892 => x"51881208",
   893 => x"52712d81",
   894 => x"f25190d6",
   895 => x"2d80d5d4",
   896 => x"08812a70",
   897 => x"81065152",
   898 => x"71a43880",
   899 => x"d4840851",
   900 => x"90d62d80",
   901 => x"d5d40881",
   902 => x"2a708106",
   903 => x"5152718e",
   904 => x"3880d6ac",
   905 => x"08820652",
   906 => x"80722580",
   907 => x"c33880d6",
   908 => x"ac088206",
   909 => x"52807225",
   910 => x"843892f1",
   911 => x"2d80d6bc",
   912 => x"08ff1180",
   913 => x"d6c00856",
   914 => x"53537372",
   915 => x"258a3881",
   916 => x"1480d6c0",
   917 => x"0c9cf004",
   918 => x"72101370",
   919 => x"84291651",
   920 => x"52881208",
   921 => x"802e8938",
   922 => x"fe518812",
   923 => x"0852712d",
   924 => x"81fd5190",
   925 => x"d62d80d5",
   926 => x"d408812a",
   927 => x"70810651",
   928 => x"5271a438",
   929 => x"80d48808",
   930 => x"5190d62d",
   931 => x"80d5d408",
   932 => x"812a7081",
   933 => x"06515271",
   934 => x"8e3880d6",
   935 => x"ac088406",
   936 => x"52807225",
   937 => x"80c03880",
   938 => x"d6ac0884",
   939 => x"06528072",
   940 => x"25843892",
   941 => x"f12d80d6",
   942 => x"c008802e",
   943 => x"8a38800b",
   944 => x"80d6c00c",
   945 => x"9de60480",
   946 => x"d6bc0810",
   947 => x"80d6bc08",
   948 => x"05708429",
   949 => x"16515288",
   950 => x"1208802e",
   951 => x"8938fd51",
   952 => x"88120852",
   953 => x"712d81fa",
   954 => x"5190d62d",
   955 => x"80d5d408",
   956 => x"812a7081",
   957 => x"06515271",
   958 => x"a43880d4",
   959 => x"8c085190",
   960 => x"d62d80d5",
   961 => x"d408812a",
   962 => x"70810651",
   963 => x"52718e38",
   964 => x"80d6ac08",
   965 => x"88065280",
   966 => x"722580c0",
   967 => x"3880d6ac",
   968 => x"08880652",
   969 => x"80722584",
   970 => x"3892f12d",
   971 => x"80d6bc08",
   972 => x"ff115452",
   973 => x"80d6c008",
   974 => x"73258938",
   975 => x"7280d6c0",
   976 => x"0c9edc04",
   977 => x"71101270",
   978 => x"84291651",
   979 => x"52881208",
   980 => x"802e8938",
   981 => x"fc518812",
   982 => x"0852712d",
   983 => x"80d6c008",
   984 => x"70535473",
   985 => x"802e8a38",
   986 => x"8c15ff15",
   987 => x"55559ee3",
   988 => x"04820b80",
   989 => x"d5e80c71",
   990 => x"8f0680d5",
   991 => x"e40c81eb",
   992 => x"5190d62d",
   993 => x"80d5d408",
   994 => x"812a7081",
   995 => x"06515271",
   996 => x"802ead38",
   997 => x"7408852e",
   998 => x"098106a4",
   999 => x"38881580",
  1000 => x"f52dff05",
  1001 => x"52718816",
  1002 => x"81b72d71",
  1003 => x"982b5271",
  1004 => x"80258838",
  1005 => x"800b8816",
  1006 => x"81b72d74",
  1007 => x"5193ef2d",
  1008 => x"81f45190",
  1009 => x"d62d80d5",
  1010 => x"d408812a",
  1011 => x"70810651",
  1012 => x"5271802e",
  1013 => x"b3387408",
  1014 => x"852e0981",
  1015 => x"06aa3888",
  1016 => x"1580f52d",
  1017 => x"81055271",
  1018 => x"881681b7",
  1019 => x"2d7181ff",
  1020 => x"068b1680",
  1021 => x"f52d5452",
  1022 => x"72722787",
  1023 => x"38728816",
  1024 => x"81b72d74",
  1025 => x"5193ef2d",
  1026 => x"80da5190",
  1027 => x"d62d80d5",
  1028 => x"d408812a",
  1029 => x"70810651",
  1030 => x"52718e38",
  1031 => x"80d6ac08",
  1032 => x"90065280",
  1033 => x"722581bc",
  1034 => x"3880d6b8",
  1035 => x"0880d6ac",
  1036 => x"08900653",
  1037 => x"53807225",
  1038 => x"843892f1",
  1039 => x"2d80d6c0",
  1040 => x"08547380",
  1041 => x"2e8a388c",
  1042 => x"13ff1555",
  1043 => x"53a0c204",
  1044 => x"72085271",
  1045 => x"822ea638",
  1046 => x"71822689",
  1047 => x"3871812e",
  1048 => x"aa38a1e4",
  1049 => x"0471832e",
  1050 => x"b4387184",
  1051 => x"2e098106",
  1052 => x"80f23888",
  1053 => x"13085195",
  1054 => x"c52da1e4",
  1055 => x"0480d6c0",
  1056 => x"08518813",
  1057 => x"0852712d",
  1058 => x"a1e40481",
  1059 => x"0b881408",
  1060 => x"2b80d3e8",
  1061 => x"083280d3",
  1062 => x"e80ca1b8",
  1063 => x"04881380",
  1064 => x"f52d8105",
  1065 => x"8b1480f5",
  1066 => x"2d535471",
  1067 => x"74248338",
  1068 => x"80547388",
  1069 => x"1481b72d",
  1070 => x"949f2da1",
  1071 => x"e4047508",
  1072 => x"802ea438",
  1073 => x"75085190",
  1074 => x"d62d80d5",
  1075 => x"d4088106",
  1076 => x"5271802e",
  1077 => x"8c3880d6",
  1078 => x"c0085184",
  1079 => x"16085271",
  1080 => x"2d881656",
  1081 => x"75d83880",
  1082 => x"54800b80",
  1083 => x"d5e80c73",
  1084 => x"8f0680d5",
  1085 => x"e40ca052",
  1086 => x"7380d6c0",
  1087 => x"082e0981",
  1088 => x"06993880",
  1089 => x"d6bc08ff",
  1090 => x"05743270",
  1091 => x"09810570",
  1092 => x"72079f2a",
  1093 => x"91713151",
  1094 => x"51535371",
  1095 => x"5183842d",
  1096 => x"8114548e",
  1097 => x"7425c238",
  1098 => x"80d49408",
  1099 => x"80d5d40c",
  1100 => x"0298050d",
  1101 => x"0402f405",
  1102 => x"0dd45281",
  1103 => x"ff720c71",
  1104 => x"085381ff",
  1105 => x"720c7288",
  1106 => x"2b83fe80",
  1107 => x"06720870",
  1108 => x"81ff0651",
  1109 => x"525381ff",
  1110 => x"720c7271",
  1111 => x"07882b72",
  1112 => x"087081ff",
  1113 => x"06515253",
  1114 => x"81ff720c",
  1115 => x"72710788",
  1116 => x"2b720870",
  1117 => x"81ff0672",
  1118 => x"0780d5d4",
  1119 => x"0c525302",
  1120 => x"8c050d04",
  1121 => x"02f4050d",
  1122 => x"74767181",
  1123 => x"ff06d40c",
  1124 => x"535380d6",
  1125 => x"c8088538",
  1126 => x"71892b52",
  1127 => x"71982ad4",
  1128 => x"0c71902a",
  1129 => x"7081ff06",
  1130 => x"d40c5171",
  1131 => x"882a7081",
  1132 => x"ff06d40c",
  1133 => x"517181ff",
  1134 => x"06d40c72",
  1135 => x"902a7081",
  1136 => x"ff06d40c",
  1137 => x"51d40870",
  1138 => x"81ff0651",
  1139 => x"5182b8bf",
  1140 => x"527081ff",
  1141 => x"2e098106",
  1142 => x"943881ff",
  1143 => x"0bd40cd4",
  1144 => x"087081ff",
  1145 => x"06ff1454",
  1146 => x"515171e5",
  1147 => x"387080d5",
  1148 => x"d40c028c",
  1149 => x"050d0402",
  1150 => x"fc050d81",
  1151 => x"c75181ff",
  1152 => x"0bd40cff",
  1153 => x"11517080",
  1154 => x"25f43802",
  1155 => x"84050d04",
  1156 => x"02f4050d",
  1157 => x"81ff0bd4",
  1158 => x"0c935380",
  1159 => x"5287fc80",
  1160 => x"c151a384",
  1161 => x"2d80d5d4",
  1162 => x"088b3881",
  1163 => x"ff0bd40c",
  1164 => x"8153a4be",
  1165 => x"04a3f72d",
  1166 => x"ff135372",
  1167 => x"de387280",
  1168 => x"d5d40c02",
  1169 => x"8c050d04",
  1170 => x"02ec050d",
  1171 => x"810b80d6",
  1172 => x"c80c8454",
  1173 => x"d008708f",
  1174 => x"2a708106",
  1175 => x"51515372",
  1176 => x"f33872d0",
  1177 => x"0ca3f72d",
  1178 => x"80cac451",
  1179 => x"87f12dd0",
  1180 => x"08708f2a",
  1181 => x"70810651",
  1182 => x"515372f3",
  1183 => x"38810bd0",
  1184 => x"0cb15380",
  1185 => x"5284d480",
  1186 => x"c051a384",
  1187 => x"2d80d5d4",
  1188 => x"08812e93",
  1189 => x"3872822e",
  1190 => x"bf38ff13",
  1191 => x"5372e438",
  1192 => x"ff145473",
  1193 => x"ffae38a3",
  1194 => x"f72d83aa",
  1195 => x"52849c80",
  1196 => x"c851a384",
  1197 => x"2d80d5d4",
  1198 => x"08812e09",
  1199 => x"81069338",
  1200 => x"a2b52d80",
  1201 => x"d5d40883",
  1202 => x"ffff0653",
  1203 => x"7283aa2e",
  1204 => x"9f38a490",
  1205 => x"2da5eb04",
  1206 => x"80cad051",
  1207 => x"87f12d80",
  1208 => x"53a7c004",
  1209 => x"80cae851",
  1210 => x"87f12d80",
  1211 => x"54a79104",
  1212 => x"81ff0bd4",
  1213 => x"0cb154a3",
  1214 => x"f72d8fcf",
  1215 => x"53805287",
  1216 => x"fc80f751",
  1217 => x"a3842d80",
  1218 => x"d5d40855",
  1219 => x"80d5d408",
  1220 => x"812e0981",
  1221 => x"069c3881",
  1222 => x"ff0bd40c",
  1223 => x"820a5284",
  1224 => x"9c80e951",
  1225 => x"a3842d80",
  1226 => x"d5d40880",
  1227 => x"2e8d38a3",
  1228 => x"f72dff13",
  1229 => x"5372c638",
  1230 => x"a7840481",
  1231 => x"ff0bd40c",
  1232 => x"80d5d408",
  1233 => x"5287fc80",
  1234 => x"fa51a384",
  1235 => x"2d80d5d4",
  1236 => x"08b23881",
  1237 => x"ff0bd40c",
  1238 => x"d4085381",
  1239 => x"ff0bd40c",
  1240 => x"81ff0bd4",
  1241 => x"0c81ff0b",
  1242 => x"d40c81ff",
  1243 => x"0bd40c72",
  1244 => x"862a7081",
  1245 => x"06765651",
  1246 => x"53729638",
  1247 => x"80d5d408",
  1248 => x"54a79104",
  1249 => x"73822efe",
  1250 => x"db38ff14",
  1251 => x"5473fee7",
  1252 => x"387380d6",
  1253 => x"c80c738b",
  1254 => x"38815287",
  1255 => x"fc80d051",
  1256 => x"a3842d81",
  1257 => x"ff0bd40c",
  1258 => x"d008708f",
  1259 => x"2a708106",
  1260 => x"51515372",
  1261 => x"f33872d0",
  1262 => x"0c81ff0b",
  1263 => x"d40c8153",
  1264 => x"7280d5d4",
  1265 => x"0c029405",
  1266 => x"0d0402e8",
  1267 => x"050d7855",
  1268 => x"805681ff",
  1269 => x"0bd40cd0",
  1270 => x"08708f2a",
  1271 => x"70810651",
  1272 => x"515372f3",
  1273 => x"3882810b",
  1274 => x"d00c81ff",
  1275 => x"0bd40c77",
  1276 => x"5287fc80",
  1277 => x"d151a384",
  1278 => x"2d80dbc6",
  1279 => x"df5480d5",
  1280 => x"d408802e",
  1281 => x"8b3880cb",
  1282 => x"885187f1",
  1283 => x"2da8e404",
  1284 => x"81ff0bd4",
  1285 => x"0cd40870",
  1286 => x"81ff0651",
  1287 => x"537281fe",
  1288 => x"2e098106",
  1289 => x"9e3880ff",
  1290 => x"53a2b52d",
  1291 => x"80d5d408",
  1292 => x"75708405",
  1293 => x"570cff13",
  1294 => x"53728025",
  1295 => x"ec388156",
  1296 => x"a8c904ff",
  1297 => x"145473c8",
  1298 => x"3881ff0b",
  1299 => x"d40c81ff",
  1300 => x"0bd40cd0",
  1301 => x"08708f2a",
  1302 => x"70810651",
  1303 => x"515372f3",
  1304 => x"3872d00c",
  1305 => x"7580d5d4",
  1306 => x"0c029805",
  1307 => x"0d0402e8",
  1308 => x"050d7779",
  1309 => x"7b585555",
  1310 => x"80537276",
  1311 => x"25a33874",
  1312 => x"70810556",
  1313 => x"80f52d74",
  1314 => x"70810556",
  1315 => x"80f52d52",
  1316 => x"5271712e",
  1317 => x"86388151",
  1318 => x"a9a30481",
  1319 => x"1353a8fa",
  1320 => x"04805170",
  1321 => x"80d5d40c",
  1322 => x"0298050d",
  1323 => x"0402ec05",
  1324 => x"0d765574",
  1325 => x"802e80c2",
  1326 => x"389a1580",
  1327 => x"e02d51b7",
  1328 => x"e82d80d5",
  1329 => x"d40880d5",
  1330 => x"d40880dc",
  1331 => x"fc0c80d5",
  1332 => x"d4085454",
  1333 => x"80dcd808",
  1334 => x"802e9a38",
  1335 => x"941580e0",
  1336 => x"2d51b7e8",
  1337 => x"2d80d5d4",
  1338 => x"08902b83",
  1339 => x"fff00a06",
  1340 => x"70750751",
  1341 => x"537280dc",
  1342 => x"fc0c80dc",
  1343 => x"fc085372",
  1344 => x"802e9d38",
  1345 => x"80dcd008",
  1346 => x"fe147129",
  1347 => x"80dce408",
  1348 => x"0580dd80",
  1349 => x"0c70842b",
  1350 => x"80dcdc0c",
  1351 => x"54aace04",
  1352 => x"80dce808",
  1353 => x"80dcfc0c",
  1354 => x"80dcec08",
  1355 => x"80dd800c",
  1356 => x"80dcd808",
  1357 => x"802e8b38",
  1358 => x"80dcd008",
  1359 => x"842b53aa",
  1360 => x"c90480dc",
  1361 => x"f008842b",
  1362 => x"537280dc",
  1363 => x"dc0c0294",
  1364 => x"050d0402",
  1365 => x"d8050d80",
  1366 => x"0b80dcd8",
  1367 => x"0c8454a4",
  1368 => x"c82d80d5",
  1369 => x"d408802e",
  1370 => x"973880d6",
  1371 => x"cc528051",
  1372 => x"a7ca2d80",
  1373 => x"d5d40880",
  1374 => x"2e8638fe",
  1375 => x"54ab8804",
  1376 => x"ff145473",
  1377 => x"8024d838",
  1378 => x"738d3880",
  1379 => x"cb985187",
  1380 => x"f12d7355",
  1381 => x"b0dd0480",
  1382 => x"56810b80",
  1383 => x"dd840c88",
  1384 => x"5380cbac",
  1385 => x"5280d782",
  1386 => x"51a8ee2d",
  1387 => x"80d5d408",
  1388 => x"762e0981",
  1389 => x"06893880",
  1390 => x"d5d40880",
  1391 => x"dd840c88",
  1392 => x"5380cbb8",
  1393 => x"5280d79e",
  1394 => x"51a8ee2d",
  1395 => x"80d5d408",
  1396 => x"893880d5",
  1397 => x"d40880dd",
  1398 => x"840c80dd",
  1399 => x"8408802e",
  1400 => x"81813880",
  1401 => x"da920b80",
  1402 => x"f52d80da",
  1403 => x"930b80f5",
  1404 => x"2d71982b",
  1405 => x"71902b07",
  1406 => x"80da940b",
  1407 => x"80f52d70",
  1408 => x"882b7207",
  1409 => x"80da950b",
  1410 => x"80f52d71",
  1411 => x"0780daca",
  1412 => x"0b80f52d",
  1413 => x"80dacb0b",
  1414 => x"80f52d71",
  1415 => x"882b0753",
  1416 => x"5f54525a",
  1417 => x"56575573",
  1418 => x"81abaa2e",
  1419 => x"0981068e",
  1420 => x"387551b7",
  1421 => x"b72d80d5",
  1422 => x"d40856ac",
  1423 => x"cc047382",
  1424 => x"d4d52e88",
  1425 => x"3880cbc4",
  1426 => x"51ad9804",
  1427 => x"80d6cc52",
  1428 => x"7551a7ca",
  1429 => x"2d80d5d4",
  1430 => x"085580d5",
  1431 => x"d408802e",
  1432 => x"83fb3888",
  1433 => x"5380cbb8",
  1434 => x"5280d79e",
  1435 => x"51a8ee2d",
  1436 => x"80d5d408",
  1437 => x"8a38810b",
  1438 => x"80dcd80c",
  1439 => x"ad9e0488",
  1440 => x"5380cbac",
  1441 => x"5280d782",
  1442 => x"51a8ee2d",
  1443 => x"80d5d408",
  1444 => x"802e8b38",
  1445 => x"80cbd851",
  1446 => x"87f12dad",
  1447 => x"fd0480da",
  1448 => x"ca0b80f5",
  1449 => x"2d547380",
  1450 => x"d52e0981",
  1451 => x"0680ce38",
  1452 => x"80dacb0b",
  1453 => x"80f52d54",
  1454 => x"7381aa2e",
  1455 => x"098106bd",
  1456 => x"38800b80",
  1457 => x"d6cc0b80",
  1458 => x"f52d5654",
  1459 => x"7481e92e",
  1460 => x"83388154",
  1461 => x"7481eb2e",
  1462 => x"8c388055",
  1463 => x"73752e09",
  1464 => x"810682f9",
  1465 => x"3880d6d7",
  1466 => x"0b80f52d",
  1467 => x"55748e38",
  1468 => x"80d6d80b",
  1469 => x"80f52d54",
  1470 => x"73822e86",
  1471 => x"388055b0",
  1472 => x"dd0480d6",
  1473 => x"d90b80f5",
  1474 => x"2d7080dc",
  1475 => x"d00cff05",
  1476 => x"80dcd40c",
  1477 => x"80d6da0b",
  1478 => x"80f52d80",
  1479 => x"d6db0b80",
  1480 => x"f52d5876",
  1481 => x"05778280",
  1482 => x"29057080",
  1483 => x"dce00c80",
  1484 => x"d6dc0b80",
  1485 => x"f52d7080",
  1486 => x"dcf40c80",
  1487 => x"dcd80859",
  1488 => x"57587680",
  1489 => x"2e81b738",
  1490 => x"885380cb",
  1491 => x"b85280d7",
  1492 => x"9e51a8ee",
  1493 => x"2d80d5d4",
  1494 => x"08828238",
  1495 => x"80dcd008",
  1496 => x"70842b80",
  1497 => x"dcdc0c70",
  1498 => x"80dcf00c",
  1499 => x"80d6f10b",
  1500 => x"80f52d80",
  1501 => x"d6f00b80",
  1502 => x"f52d7182",
  1503 => x"80290580",
  1504 => x"d6f20b80",
  1505 => x"f52d7084",
  1506 => x"80802912",
  1507 => x"80d6f30b",
  1508 => x"80f52d70",
  1509 => x"81800a29",
  1510 => x"127080dc",
  1511 => x"f80c80dc",
  1512 => x"f4087129",
  1513 => x"80dce008",
  1514 => x"057080dc",
  1515 => x"e40c80d6",
  1516 => x"f90b80f5",
  1517 => x"2d80d6f8",
  1518 => x"0b80f52d",
  1519 => x"71828029",
  1520 => x"0580d6fa",
  1521 => x"0b80f52d",
  1522 => x"70848080",
  1523 => x"291280d6",
  1524 => x"fb0b80f5",
  1525 => x"2d70982b",
  1526 => x"81f00a06",
  1527 => x"72057080",
  1528 => x"dce80cfe",
  1529 => x"117e2977",
  1530 => x"0580dcec",
  1531 => x"0c525952",
  1532 => x"43545e51",
  1533 => x"5259525d",
  1534 => x"575957b0",
  1535 => x"d60480d6",
  1536 => x"de0b80f5",
  1537 => x"2d80d6dd",
  1538 => x"0b80f52d",
  1539 => x"71828029",
  1540 => x"057080dc",
  1541 => x"dc0c70a0",
  1542 => x"2983ff05",
  1543 => x"70892a70",
  1544 => x"80dcf00c",
  1545 => x"80d6e30b",
  1546 => x"80f52d80",
  1547 => x"d6e20b80",
  1548 => x"f52d7182",
  1549 => x"80290570",
  1550 => x"80dcf80c",
  1551 => x"7b71291e",
  1552 => x"7080dcec",
  1553 => x"0c7d80dc",
  1554 => x"e80c7305",
  1555 => x"80dce40c",
  1556 => x"555e5151",
  1557 => x"55558051",
  1558 => x"a9ad2d81",
  1559 => x"557480d5",
  1560 => x"d40c02a8",
  1561 => x"050d0402",
  1562 => x"ec050d76",
  1563 => x"70872c71",
  1564 => x"80ff0655",
  1565 => x"565480dc",
  1566 => x"d8088a38",
  1567 => x"73882c74",
  1568 => x"81ff0654",
  1569 => x"5580d6cc",
  1570 => x"5280dce0",
  1571 => x"081551a7",
  1572 => x"ca2d80d5",
  1573 => x"d4085480",
  1574 => x"d5d40880",
  1575 => x"2eb83880",
  1576 => x"dcd80880",
  1577 => x"2e9a3872",
  1578 => x"842980d6",
  1579 => x"cc057008",
  1580 => x"5253b7b7",
  1581 => x"2d80d5d4",
  1582 => x"08f00a06",
  1583 => x"53b1d404",
  1584 => x"721080d6",
  1585 => x"cc057080",
  1586 => x"e02d5253",
  1587 => x"b7e82d80",
  1588 => x"d5d40853",
  1589 => x"72547380",
  1590 => x"d5d40c02",
  1591 => x"94050d04",
  1592 => x"02e0050d",
  1593 => x"7970842c",
  1594 => x"80dd8008",
  1595 => x"05718f06",
  1596 => x"52555372",
  1597 => x"8a3880d6",
  1598 => x"cc527351",
  1599 => x"a7ca2d72",
  1600 => x"a02980d6",
  1601 => x"cc055480",
  1602 => x"7480f52d",
  1603 => x"56537473",
  1604 => x"2e833881",
  1605 => x"537481e5",
  1606 => x"2e81f438",
  1607 => x"81707406",
  1608 => x"54587280",
  1609 => x"2e81e838",
  1610 => x"8b1480f5",
  1611 => x"2d70832a",
  1612 => x"79065856",
  1613 => x"769b3880",
  1614 => x"d4980853",
  1615 => x"72893872",
  1616 => x"80dacc0b",
  1617 => x"81b72d76",
  1618 => x"80d4980c",
  1619 => x"7353b491",
  1620 => x"04758f2e",
  1621 => x"09810681",
  1622 => x"b638749f",
  1623 => x"068d2980",
  1624 => x"dabf1151",
  1625 => x"53811480",
  1626 => x"f52d7370",
  1627 => x"81055581",
  1628 => x"b72d8314",
  1629 => x"80f52d73",
  1630 => x"70810555",
  1631 => x"81b72d85",
  1632 => x"1480f52d",
  1633 => x"73708105",
  1634 => x"5581b72d",
  1635 => x"871480f5",
  1636 => x"2d737081",
  1637 => x"055581b7",
  1638 => x"2d891480",
  1639 => x"f52d7370",
  1640 => x"81055581",
  1641 => x"b72d8e14",
  1642 => x"80f52d73",
  1643 => x"70810555",
  1644 => x"81b72d90",
  1645 => x"1480f52d",
  1646 => x"73708105",
  1647 => x"5581b72d",
  1648 => x"921480f5",
  1649 => x"2d737081",
  1650 => x"055581b7",
  1651 => x"2d941480",
  1652 => x"f52d7370",
  1653 => x"81055581",
  1654 => x"b72d9614",
  1655 => x"80f52d73",
  1656 => x"70810555",
  1657 => x"81b72d98",
  1658 => x"1480f52d",
  1659 => x"73708105",
  1660 => x"5581b72d",
  1661 => x"9c1480f5",
  1662 => x"2d737081",
  1663 => x"055581b7",
  1664 => x"2d9e1480",
  1665 => x"f52d7381",
  1666 => x"b72d7780",
  1667 => x"d4980c80",
  1668 => x"537280d5",
  1669 => x"d40c02a0",
  1670 => x"050d0402",
  1671 => x"cc050d7e",
  1672 => x"605e5b80",
  1673 => x"0b80dcfc",
  1674 => x"0880dd80",
  1675 => x"08595d56",
  1676 => x"805980dc",
  1677 => x"dc08792e",
  1678 => x"81de3878",
  1679 => x"8f06a017",
  1680 => x"57547391",
  1681 => x"3880d6cc",
  1682 => x"52765181",
  1683 => x"1757a7ca",
  1684 => x"2d80d6cc",
  1685 => x"56807680",
  1686 => x"f52d5654",
  1687 => x"74742e83",
  1688 => x"38815474",
  1689 => x"81e52e81",
  1690 => x"a3388170",
  1691 => x"7506555a",
  1692 => x"73802e81",
  1693 => x"97388b16",
  1694 => x"80f52d70",
  1695 => x"98065954",
  1696 => x"7780e338",
  1697 => x"8b537c52",
  1698 => x"7551a8ee",
  1699 => x"2d80d5d4",
  1700 => x"0880f938",
  1701 => x"9c160851",
  1702 => x"b7b72d80",
  1703 => x"d5d40884",
  1704 => x"1c0c9a16",
  1705 => x"80e02d51",
  1706 => x"b7e82d80",
  1707 => x"d5d40880",
  1708 => x"d5d40888",
  1709 => x"1d0c80d5",
  1710 => x"d4085555",
  1711 => x"80dcd808",
  1712 => x"802e9938",
  1713 => x"941680e0",
  1714 => x"2d51b7e8",
  1715 => x"2d80d5d4",
  1716 => x"08902b83",
  1717 => x"fff00a06",
  1718 => x"70165154",
  1719 => x"73881c0c",
  1720 => x"777b0cb6",
  1721 => x"87047384",
  1722 => x"2a708106",
  1723 => x"51547380",
  1724 => x"2e9a388b",
  1725 => x"537c5275",
  1726 => x"51a8ee2d",
  1727 => x"80d5d408",
  1728 => x"8b387551",
  1729 => x"a9ad2d79",
  1730 => x"54b6d404",
  1731 => x"81195980",
  1732 => x"dcdc0879",
  1733 => x"26fea438",
  1734 => x"80dcd808",
  1735 => x"802eb338",
  1736 => x"7b51b0e7",
  1737 => x"2d80d5d4",
  1738 => x"0880d5d4",
  1739 => x"0880ffff",
  1740 => x"fff80655",
  1741 => x"5c7380ff",
  1742 => x"fffff82e",
  1743 => x"953880d5",
  1744 => x"d408fe05",
  1745 => x"80dcd008",
  1746 => x"2980dce4",
  1747 => x"080557b4",
  1748 => x"b0048054",
  1749 => x"7380d5d4",
  1750 => x"0c02b405",
  1751 => x"0d0402f4",
  1752 => x"050d7470",
  1753 => x"08810571",
  1754 => x"0c700880",
  1755 => x"dcd40806",
  1756 => x"5353718f",
  1757 => x"38881308",
  1758 => x"51b0e72d",
  1759 => x"80d5d408",
  1760 => x"88140c81",
  1761 => x"0b80d5d4",
  1762 => x"0c028c05",
  1763 => x"0d0402f0",
  1764 => x"050d7588",
  1765 => x"1108fe05",
  1766 => x"80dcd008",
  1767 => x"2980dce4",
  1768 => x"08117208",
  1769 => x"80dcd408",
  1770 => x"06057955",
  1771 => x"535454a7",
  1772 => x"ca2d0290",
  1773 => x"050d0402",
  1774 => x"f4050d74",
  1775 => x"70882a83",
  1776 => x"fe800670",
  1777 => x"72982a07",
  1778 => x"72882b87",
  1779 => x"fc808006",
  1780 => x"73982b81",
  1781 => x"f00a0671",
  1782 => x"73070780",
  1783 => x"d5d40c56",
  1784 => x"51535102",
  1785 => x"8c050d04",
  1786 => x"02f8050d",
  1787 => x"028e0580",
  1788 => x"f52d7488",
  1789 => x"2b077083",
  1790 => x"ffff0680",
  1791 => x"d5d40c51",
  1792 => x"0288050d",
  1793 => x"0402ec05",
  1794 => x"0d76787a",
  1795 => x"53555381",
  1796 => x"55807125",
  1797 => x"ae387052",
  1798 => x"73708105",
  1799 => x"5580f52d",
  1800 => x"73708105",
  1801 => x"5581b72d",
  1802 => x"7380f52d",
  1803 => x"51708638",
  1804 => x"7055b8b8",
  1805 => x"04748638",
  1806 => x"a07381b7",
  1807 => x"2dff1252",
  1808 => x"71d63880",
  1809 => x"7381b72d",
  1810 => x"0294050d",
  1811 => x"0402e805",
  1812 => x"0d775680",
  1813 => x"70565473",
  1814 => x"7624b638",
  1815 => x"80dcdc08",
  1816 => x"742eae38",
  1817 => x"7351b1e0",
  1818 => x"2d80d5d4",
  1819 => x"0880d5d4",
  1820 => x"08098105",
  1821 => x"7080d5d4",
  1822 => x"08079f2a",
  1823 => x"77058117",
  1824 => x"57575353",
  1825 => x"74762489",
  1826 => x"3880dcdc",
  1827 => x"087426d4",
  1828 => x"387280d5",
  1829 => x"d40c0298",
  1830 => x"050d0402",
  1831 => x"f0050d80",
  1832 => x"d5d00816",
  1833 => x"51b8cd2d",
  1834 => x"80d5d408",
  1835 => x"802e9f38",
  1836 => x"8b5380d5",
  1837 => x"d4085280",
  1838 => x"dacc51b8",
  1839 => x"852d80dd",
  1840 => x"88085473",
  1841 => x"802e8738",
  1842 => x"80dacc51",
  1843 => x"732d0290",
  1844 => x"050d0402",
  1845 => x"dc050d80",
  1846 => x"705a5574",
  1847 => x"80d5d008",
  1848 => x"25b43880",
  1849 => x"dcdc0875",
  1850 => x"2eac3878",
  1851 => x"51b1e02d",
  1852 => x"80d5d408",
  1853 => x"09810570",
  1854 => x"80d5d408",
  1855 => x"079f2a76",
  1856 => x"05811b5b",
  1857 => x"56547480",
  1858 => x"d5d00825",
  1859 => x"893880dc",
  1860 => x"dc087926",
  1861 => x"d6388055",
  1862 => x"7880dcdc",
  1863 => x"082781db",
  1864 => x"387851b1",
  1865 => x"e02d80d5",
  1866 => x"d408802e",
  1867 => x"81ad3880",
  1868 => x"d5d4088b",
  1869 => x"0580f52d",
  1870 => x"70842a70",
  1871 => x"81067710",
  1872 => x"78842b80",
  1873 => x"dacc0b80",
  1874 => x"f52d5c5c",
  1875 => x"53515556",
  1876 => x"73802e80",
  1877 => x"cb387416",
  1878 => x"822bbc9f",
  1879 => x"0b80d4a4",
  1880 => x"120c5477",
  1881 => x"75311080",
  1882 => x"dd8c1155",
  1883 => x"56907470",
  1884 => x"81055681",
  1885 => x"b72da074",
  1886 => x"81b72d76",
  1887 => x"81ff0681",
  1888 => x"16585473",
  1889 => x"802e8a38",
  1890 => x"9c5380da",
  1891 => x"cc52bb98",
  1892 => x"048b5380",
  1893 => x"d5d40852",
  1894 => x"80dd8e16",
  1895 => x"51bbd304",
  1896 => x"7416822b",
  1897 => x"b99b0b80",
  1898 => x"d4a4120c",
  1899 => x"547681ff",
  1900 => x"06811658",
  1901 => x"5473802e",
  1902 => x"8a389c53",
  1903 => x"80dacc52",
  1904 => x"bbca048b",
  1905 => x"5380d5d4",
  1906 => x"08527775",
  1907 => x"311080dd",
  1908 => x"8c055176",
  1909 => x"55b8852d",
  1910 => x"bbf00474",
  1911 => x"90297531",
  1912 => x"701080dd",
  1913 => x"8c055154",
  1914 => x"80d5d408",
  1915 => x"7481b72d",
  1916 => x"81195974",
  1917 => x"8b24a338",
  1918 => x"ba980474",
  1919 => x"90297531",
  1920 => x"701080dd",
  1921 => x"8c058c77",
  1922 => x"31575154",
  1923 => x"807481b7",
  1924 => x"2d9e14ff",
  1925 => x"16565474",
  1926 => x"f33802a4",
  1927 => x"050d0402",
  1928 => x"fc050d80",
  1929 => x"d5d00813",
  1930 => x"51b8cd2d",
  1931 => x"80d5d408",
  1932 => x"802e8938",
  1933 => x"80d5d408",
  1934 => x"51a9ad2d",
  1935 => x"800b80d5",
  1936 => x"d00cb9d3",
  1937 => x"2d949f2d",
  1938 => x"0284050d",
  1939 => x"0402f805",
  1940 => x"0d735170",
  1941 => x"fd2eb138",
  1942 => x"70fd248a",
  1943 => x"3870fc2e",
  1944 => x"80cd38bd",
  1945 => x"c90470fe",
  1946 => x"2eb83870",
  1947 => x"ff2e0981",
  1948 => x"0680d638",
  1949 => x"80d5d008",
  1950 => x"5170802e",
  1951 => x"80cb38ff",
  1952 => x"1180d5d0",
  1953 => x"0cbdc904",
  1954 => x"80d5d008",
  1955 => x"f4057080",
  1956 => x"d5d00c51",
  1957 => x"708025b1",
  1958 => x"38800b80",
  1959 => x"d5d00cbd",
  1960 => x"c90480d5",
  1961 => x"d0088105",
  1962 => x"80d5d00c",
  1963 => x"bdc90480",
  1964 => x"d5d0088c",
  1965 => x"117080d5",
  1966 => x"d00c5252",
  1967 => x"80dcdc08",
  1968 => x"71268638",
  1969 => x"7180d5d0",
  1970 => x"0cb9d32d",
  1971 => x"949f2d02",
  1972 => x"88050d04",
  1973 => x"02fc050d",
  1974 => x"800b80d5",
  1975 => x"d00cb9d3",
  1976 => x"2d93882d",
  1977 => x"80d5d408",
  1978 => x"80d5c00c",
  1979 => x"80d49c51",
  1980 => x"95c52d02",
  1981 => x"84050d04",
  1982 => x"02f8050d",
  1983 => x"810b80cd",
  1984 => x"e40c80d5",
  1985 => x"fc08bff9",
  1986 => x"ff068180",
  1987 => x"077080d5",
  1988 => x"fc0cfc0c",
  1989 => x"7351bdd4",
  1990 => x"2d028805",
  1991 => x"0d0402f8",
  1992 => x"050d820b",
  1993 => x"80cde40c",
  1994 => x"80d5fc08",
  1995 => x"bffaff06",
  1996 => x"82800770",
  1997 => x"80d5fc0c",
  1998 => x"fc0c7351",
  1999 => x"bdd42d02",
  2000 => x"88050d04",
  2001 => x"02f8050d",
  2002 => x"830b80cd",
  2003 => x"e40c80d5",
  2004 => x"fc08bfff",
  2005 => x"ff068780",
  2006 => x"077080d5",
  2007 => x"fc0cfc0c",
  2008 => x"7351bdd4",
  2009 => x"2d028805",
  2010 => x"0d047180",
  2011 => x"dd880c04",
  2012 => x"00ffffff",
  2013 => x"ff00ffff",
  2014 => x"ffff00ff",
  2015 => x"ffffff00",
  2016 => x"54686572",
  2017 => x"65206973",
  2018 => x"206e6f20",
  2019 => x"696d6167",
  2020 => x"65207768",
  2021 => x"656e206c",
  2022 => x"6f616469",
  2023 => x"6e670000",
  2024 => x"436f6e74",
  2025 => x"696e7565",
  2026 => x"00000000",
  2027 => x"3d205a58",
  2028 => x"38312f5a",
  2029 => x"58383020",
  2030 => x"436f6e66",
  2031 => x"69677572",
  2032 => x"6174696f",
  2033 => x"6e203d00",
  2034 => x"3d3d3d3d",
  2035 => x"3d3d3d3d",
  2036 => x"3d3d3d3d",
  2037 => x"3d3d3d3d",
  2038 => x"3d3d3d3d",
  2039 => x"3d3d3d3d",
  2040 => x"3d3d3d00",
  2041 => x"4c6f7720",
  2042 => x"52414d3a",
  2043 => x"204f6666",
  2044 => x"2f384b42",
  2045 => x"00000000",
  2046 => x"51532043",
  2047 => x"4852533a",
  2048 => x"44697361",
  2049 => x"626c6564",
  2050 => x"2f456e61",
  2051 => x"626c6564",
  2052 => x"28463129",
  2053 => x"00000000",
  2054 => x"4348524f",
  2055 => x"4d413831",
  2056 => x"3a204469",
  2057 => x"7361626c",
  2058 => x"65642f45",
  2059 => x"6e61626c",
  2060 => x"65640000",
  2061 => x"496e7665",
  2062 => x"72736520",
  2063 => x"76696465",
  2064 => x"6f3a204f",
  2065 => x"66662f4f",
  2066 => x"6e000000",
  2067 => x"426c6163",
  2068 => x"6b20626f",
  2069 => x"72646572",
  2070 => x"3a204f66",
  2071 => x"662f4f6e",
  2072 => x"00000000",
  2073 => x"56696465",
  2074 => x"6f206672",
  2075 => x"65717565",
  2076 => x"6e63793a",
  2077 => x"20353048",
  2078 => x"7a2f3630",
  2079 => x"487a0000",
  2080 => x"476f2042",
  2081 => x"61636b00",
  2082 => x"536c6f77",
  2083 => x"206d6f64",
  2084 => x"65207370",
  2085 => x"6565643a",
  2086 => x"204f7269",
  2087 => x"67696e61",
  2088 => x"6c000000",
  2089 => x"536c6f77",
  2090 => x"206d6f64",
  2091 => x"65207370",
  2092 => x"6565643a",
  2093 => x"204e6f57",
  2094 => x"61697400",
  2095 => x"536c6f77",
  2096 => x"206d6f64",
  2097 => x"65207370",
  2098 => x"6565643a",
  2099 => x"20783200",
  2100 => x"536c6f77",
  2101 => x"206d6f64",
  2102 => x"65207370",
  2103 => x"6565643a",
  2104 => x"20783800",
  2105 => x"43485224",
  2106 => x"3132382f",
  2107 => x"5544473a",
  2108 => x"20313238",
  2109 => x"20436861",
  2110 => x"72730000",
  2111 => x"43485224",
  2112 => x"3132382f",
  2113 => x"5544473a",
  2114 => x"20363420",
  2115 => x"43686172",
  2116 => x"73000000",
  2117 => x"43485224",
  2118 => x"3132382f",
  2119 => x"5544473a",
  2120 => x"20446973",
  2121 => x"61626c65",
  2122 => x"64000000",
  2123 => x"4a6f7973",
  2124 => x"7469636b",
  2125 => x"3a204375",
  2126 => x"72736f72",
  2127 => x"00000000",
  2128 => x"4a6f7973",
  2129 => x"7469636b",
  2130 => x"3a205369",
  2131 => x"6e636c61",
  2132 => x"69720000",
  2133 => x"4a6f7973",
  2134 => x"7469636b",
  2135 => x"3a205a58",
  2136 => x"38310000",
  2137 => x"4d61696e",
  2138 => x"2052414d",
  2139 => x"3a203136",
  2140 => x"4b420000",
  2141 => x"4d61696e",
  2142 => x"2052414d",
  2143 => x"3a203332",
  2144 => x"4b420000",
  2145 => x"4d61696e",
  2146 => x"2052414d",
  2147 => x"3a203438",
  2148 => x"4b420000",
  2149 => x"4d61696e",
  2150 => x"2052414d",
  2151 => x"3a20314b",
  2152 => x"42000000",
  2153 => x"436f6d70",
  2154 => x"75746572",
  2155 => x"204d6f64",
  2156 => x"656c3a20",
  2157 => x"5a583831",
  2158 => x"00000000",
  2159 => x"436f6d70",
  2160 => x"75746572",
  2161 => x"204d6f64",
  2162 => x"656c3a20",
  2163 => x"5a583830",
  2164 => x"00000000",
  2165 => x"3d3d205a",
  2166 => x"5838312f",
  2167 => x"5a583830",
  2168 => x"20666f72",
  2169 => x"205a5844",
  2170 => x"4f53203d",
  2171 => x"3d000000",
  2172 => x"3d3d3d3d",
  2173 => x"3d3d3d3d",
  2174 => x"3d3d3d3d",
  2175 => x"3d3d3d3d",
  2176 => x"3d3d3d3d",
  2177 => x"3d3d3d3d",
  2178 => x"3d000000",
  2179 => x"52657365",
  2180 => x"74000000",
  2181 => x"4c6f6164",
  2182 => x"20546170",
  2183 => x"6520282e",
  2184 => x"70292010",
  2185 => x"00000000",
  2186 => x"4c6f6164",
  2187 => x"20546170",
  2188 => x"6520282e",
  2189 => x"6f292010",
  2190 => x"00000000",
  2191 => x"4c6f6164",
  2192 => x"20526f6d",
  2193 => x"2020282e",
  2194 => x"726f6d29",
  2195 => x"20100000",
  2196 => x"436f6e66",
  2197 => x"69677572",
  2198 => x"6174696f",
  2199 => x"6e206f70",
  2200 => x"74696f6e",
  2201 => x"73201000",
  2202 => x"4b657962",
  2203 => x"6f617264",
  2204 => x"2048656c",
  2205 => x"70000000",
  2206 => x"45786974",
  2207 => x"00000000",
  2208 => x"3d3d205a",
  2209 => x"5838312f",
  2210 => x"5a583830",
  2211 => x"20666f72",
  2212 => x"205a5855",
  2213 => x"4e4f203d",
  2214 => x"3d000000",
  2215 => x"524f4d20",
  2216 => x"6c6f6164",
  2217 => x"696e6720",
  2218 => x"6661696c",
  2219 => x"65640000",
  2220 => x"4f4b0000",
  2221 => x"54617065",
  2222 => x"2066696c",
  2223 => x"65204c6f",
  2224 => x"61646564",
  2225 => x"2e000000",
  2226 => x"54797065",
  2227 => x"204c4f41",
  2228 => x"44202222",
  2229 => x"202b2045",
  2230 => x"4e544552",
  2231 => x"206f6e20",
  2232 => x"5a583831",
  2233 => x"00000000",
  2234 => x"3d205a58",
  2235 => x"38312f5a",
  2236 => x"58383020",
  2237 => x"4b657962",
  2238 => x"6f617264",
  2239 => x"2048656c",
  2240 => x"70203d00",
  2241 => x"5363726f",
  2242 => x"6c6c204c",
  2243 => x"6f636b3a",
  2244 => x"20636861",
  2245 => x"6e676520",
  2246 => x"62657477",
  2247 => x"65656e00",
  2248 => x"52474220",
  2249 => x"616e6420",
  2250 => x"56474120",
  2251 => x"76696465",
  2252 => x"6f206d6f",
  2253 => x"64650000",
  2254 => x"4374726c",
  2255 => x"2b416c74",
  2256 => x"2b44656c",
  2257 => x"6574653a",
  2258 => x"20536f66",
  2259 => x"74205265",
  2260 => x"73657400",
  2261 => x"4374726c",
  2262 => x"2b416c74",
  2263 => x"2b426163",
  2264 => x"6b737061",
  2265 => x"63653a20",
  2266 => x"48617264",
  2267 => x"20726573",
  2268 => x"65740000",
  2269 => x"45736320",
  2270 => x"6f72206a",
  2271 => x"6f797374",
  2272 => x"69636b20",
  2273 => x"62742e32",
  2274 => x"3a20746f",
  2275 => x"2073686f",
  2276 => x"77000000",
  2277 => x"6f722068",
  2278 => x"69646520",
  2279 => x"74686520",
  2280 => x"6f707469",
  2281 => x"6f6e7320",
  2282 => x"6d656e75",
  2283 => x"2e000000",
  2284 => x"57415344",
  2285 => x"202f2063",
  2286 => x"7572736f",
  2287 => x"72206b65",
  2288 => x"7973202f",
  2289 => x"206a6f79",
  2290 => x"73746963",
  2291 => x"6b000000",
  2292 => x"746f2073",
  2293 => x"656c6563",
  2294 => x"74206d65",
  2295 => x"6e75206f",
  2296 => x"7074696f",
  2297 => x"6e2e0000",
  2298 => x"456e7465",
  2299 => x"72202f20",
  2300 => x"46697265",
  2301 => x"20746f20",
  2302 => x"63686f6f",
  2303 => x"7365206f",
  2304 => x"7074696f",
  2305 => x"6e2e0000",
  2306 => x"3d205a58",
  2307 => x"38312f5a",
  2308 => x"58383020",
  2309 => x"436f7265",
  2310 => x"20437265",
  2311 => x"64697473",
  2312 => x"20203d00",
  2313 => x"5a583831",
  2314 => x"2f5a5838",
  2315 => x"3020636f",
  2316 => x"72652066",
  2317 => x"6f72205a",
  2318 => x"58554e4f",
  2319 => x"2c200000",
  2320 => x"5a58444f",
  2321 => x"5320616e",
  2322 => x"64205a58",
  2323 => x"444f532b",
  2324 => x"20626f61",
  2325 => x"7264732e",
  2326 => x"00000000",
  2327 => x"4f726967",
  2328 => x"696e616c",
  2329 => x"20636f72",
  2330 => x"65732062",
  2331 => x"793a0000",
  2332 => x"202d2053",
  2333 => x"7a6f6d62",
  2334 => x"61746865",
  2335 => x"6c796920",
  2336 => x"47796f72",
  2337 => x"67792028",
  2338 => x"4d697374",
  2339 => x"29000000",
  2340 => x"202d2053",
  2341 => x"6f726765",
  2342 => x"6c696720",
  2343 => x"284d6973",
  2344 => x"74657229",
  2345 => x"00000000",
  2346 => x"506f7274",
  2347 => x"206d6164",
  2348 => x"65206279",
  2349 => x"3a204176",
  2350 => x"6c697841",
  2351 => x"00000000",
  2352 => x"496e6974",
  2353 => x"69616c69",
  2354 => x"7a696e67",
  2355 => x"20534420",
  2356 => x"63617264",
  2357 => x"0a000000",
  2358 => x"4c6f6164",
  2359 => x"696e6720",
  2360 => x"696e6974",
  2361 => x"69616c20",
  2362 => x"524f4d2e",
  2363 => x"2e2e0a00",
  2364 => x"5a583831",
  2365 => x"20202020",
  2366 => x"20202000",
  2367 => x"524f4d53",
  2368 => x"20202020",
  2369 => x"20202000",
  2370 => x"5a583858",
  2371 => x"20202020",
  2372 => x"524f4d00",
  2373 => x"4572726f",
  2374 => x"72204c6f",
  2375 => x"6164696e",
  2376 => x"6720524f",
  2377 => x"4d2e2e2e",
  2378 => x"0a000000",
  2379 => x"2e2e2020",
  2380 => x"20202020",
  2381 => x"20202000",
  2382 => x"16200000",
  2383 => x"14200000",
  2384 => x"15200000",
  2385 => x"53442069",
  2386 => x"6e69742e",
  2387 => x"2e2e0a00",
  2388 => x"53442063",
  2389 => x"61726420",
  2390 => x"72657365",
  2391 => x"74206661",
  2392 => x"696c6564",
  2393 => x"210a0000",
  2394 => x"53444843",
  2395 => x"20657272",
  2396 => x"6f72210a",
  2397 => x"00000000",
  2398 => x"57726974",
  2399 => x"65206661",
  2400 => x"696c6564",
  2401 => x"0a000000",
  2402 => x"52656164",
  2403 => x"20666169",
  2404 => x"6c65640a",
  2405 => x"00000000",
  2406 => x"43617264",
  2407 => x"20696e69",
  2408 => x"74206661",
  2409 => x"696c6564",
  2410 => x"0a000000",
  2411 => x"46415431",
  2412 => x"36202020",
  2413 => x"00000000",
  2414 => x"46415433",
  2415 => x"32202020",
  2416 => x"00000000",
  2417 => x"4e6f2070",
  2418 => x"61727469",
  2419 => x"74696f6e",
  2420 => x"20736967",
  2421 => x"0a000000",
  2422 => x"42616420",
  2423 => x"70617274",
  2424 => x"0a000000",
  2425 => x"4261636b",
  2426 => x"00000000",
  2427 => x"00000002",
  2428 => x"00000002",
  2429 => x"00001fac",
  2430 => x"00000342",
  2431 => x"00000002",
  2432 => x"00001fc8",
  2433 => x"00000342",
  2434 => x"00000003",
  2435 => x"000026dc",
  2436 => x"00000002",
  2437 => x"00000003",
  2438 => x"000026cc",
  2439 => x"00000004",
  2440 => x"00000001",
  2441 => x"00001fe4",
  2442 => x"00000000",
  2443 => x"00000003",
  2444 => x"000026c0",
  2445 => x"00000003",
  2446 => x"00000001",
  2447 => x"00001ff8",
  2448 => x"00000001",
  2449 => x"00000003",
  2450 => x"000026b4",
  2451 => x"00000003",
  2452 => x"00000001",
  2453 => x"00002018",
  2454 => x"00000002",
  2455 => x"00000001",
  2456 => x"00002034",
  2457 => x"00000003",
  2458 => x"00000001",
  2459 => x"0000204c",
  2460 => x"00000004",
  2461 => x"00000003",
  2462 => x"000026a4",
  2463 => x"00000003",
  2464 => x"00000001",
  2465 => x"00002064",
  2466 => x"00000005",
  2467 => x"00000004",
  2468 => x"00002080",
  2469 => x"00002b00",
  2470 => x"00000000",
  2471 => x"00000000",
  2472 => x"00000000",
  2473 => x"00002088",
  2474 => x"000020a4",
  2475 => x"000020bc",
  2476 => x"000020d0",
  2477 => x"000020e4",
  2478 => x"000020fc",
  2479 => x"00002114",
  2480 => x"0000212c",
  2481 => x"00002140",
  2482 => x"00002154",
  2483 => x"00002164",
  2484 => x"00002174",
  2485 => x"00002184",
  2486 => x"00002194",
  2487 => x"000021a4",
  2488 => x"000021bc",
  2489 => x"00000000",
  2490 => x"00000002",
  2491 => x"000021d4",
  2492 => x"00000343",
  2493 => x"00000002",
  2494 => x"000021f0",
  2495 => x"00000343",
  2496 => x"00000002",
  2497 => x"0000220c",
  2498 => x"00000386",
  2499 => x"00000002",
  2500 => x"00002214",
  2501 => x"00001ef8",
  2502 => x"00000002",
  2503 => x"00002228",
  2504 => x"00001f1e",
  2505 => x"00000002",
  2506 => x"0000223c",
  2507 => x"00001f44",
  2508 => x"00000002",
  2509 => x"00002250",
  2510 => x"00000353",
  2511 => x"00000002",
  2512 => x"00002268",
  2513 => x"00000363",
  2514 => x"00000002",
  2515 => x"00002278",
  2516 => x"000009a5",
  2517 => x"00000000",
  2518 => x"00000000",
  2519 => x"00000000",
  2520 => x"00000002",
  2521 => x"00002280",
  2522 => x"00000343",
  2523 => x"00000002",
  2524 => x"000021f0",
  2525 => x"00000343",
  2526 => x"00000002",
  2527 => x"0000220c",
  2528 => x"00000386",
  2529 => x"00000002",
  2530 => x"00002214",
  2531 => x"00001ef8",
  2532 => x"00000002",
  2533 => x"00002228",
  2534 => x"00001f1e",
  2535 => x"00000002",
  2536 => x"0000223c",
  2537 => x"00001f44",
  2538 => x"00000002",
  2539 => x"00002250",
  2540 => x"00000353",
  2541 => x"00000002",
  2542 => x"00002268",
  2543 => x"00000363",
  2544 => x"00000002",
  2545 => x"00002278",
  2546 => x"000009a5",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00000004",
  2551 => x"0000229c",
  2552 => x"000027d8",
  2553 => x"00000004",
  2554 => x"000022b0",
  2555 => x"00002b00",
  2556 => x"00000000",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000004",
  2560 => x"000022b4",
  2561 => x"000027fc",
  2562 => x"00000004",
  2563 => x"000022c8",
  2564 => x"000027fc",
  2565 => x"00000004",
  2566 => x"00002574",
  2567 => x"000027fc",
  2568 => x"00000004",
  2569 => x"00001f80",
  2570 => x"000027fc",
  2571 => x"00000004",
  2572 => x"00002574",
  2573 => x"000027fc",
  2574 => x"00000004",
  2575 => x"00001fa0",
  2576 => x"00002b00",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000002",
  2581 => x"000022e8",
  2582 => x"00000342",
  2583 => x"00000002",
  2584 => x"00001fc8",
  2585 => x"00000342",
  2586 => x"00000002",
  2587 => x"00002304",
  2588 => x"00000342",
  2589 => x"00000002",
  2590 => x"00002320",
  2591 => x"00000342",
  2592 => x"00000002",
  2593 => x"00002338",
  2594 => x"00000342",
  2595 => x"00000002",
  2596 => x"00002354",
  2597 => x"00000342",
  2598 => x"00000002",
  2599 => x"00002374",
  2600 => x"00000342",
  2601 => x"00000002",
  2602 => x"00002394",
  2603 => x"00000342",
  2604 => x"00000002",
  2605 => x"000023b0",
  2606 => x"00000342",
  2607 => x"00000002",
  2608 => x"000023d0",
  2609 => x"00000342",
  2610 => x"00000002",
  2611 => x"000023e8",
  2612 => x"00000342",
  2613 => x"00000002",
  2614 => x"00002574",
  2615 => x"00000342",
  2616 => x"00000004",
  2617 => x"000022b0",
  2618 => x"00002b00",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000002",
  2623 => x"00002408",
  2624 => x"00000342",
  2625 => x"00000002",
  2626 => x"00001fc8",
  2627 => x"00000342",
  2628 => x"00000002",
  2629 => x"00002424",
  2630 => x"00000342",
  2631 => x"00000002",
  2632 => x"00002440",
  2633 => x"00000342",
  2634 => x"00000002",
  2635 => x"00002574",
  2636 => x"00000342",
  2637 => x"00000002",
  2638 => x"0000245c",
  2639 => x"00000342",
  2640 => x"00000002",
  2641 => x"00002470",
  2642 => x"00000342",
  2643 => x"00000002",
  2644 => x"00002490",
  2645 => x"00000342",
  2646 => x"00000002",
  2647 => x"00002574",
  2648 => x"00000342",
  2649 => x"00000002",
  2650 => x"000024a8",
  2651 => x"00000342",
  2652 => x"00000002",
  2653 => x"00002574",
  2654 => x"00000342",
  2655 => x"00000002",
  2656 => x"00002574",
  2657 => x"00000342",
  2658 => x"00000004",
  2659 => x"000022b0",
  2660 => x"00002b00",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000006",
  2683 => x"00000043",
  2684 => x"00000042",
  2685 => x"0000003b",
  2686 => x"0000004b",
  2687 => x"0000007e",
  2688 => x"00000003",
  2689 => x"0000000b",
  2690 => x"00000083",
  2691 => x"00000023",
  2692 => x"0000007e",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000002",
  2696 => x"00002e8c",
  2697 => x"00001c9b",
  2698 => x"00000002",
  2699 => x"00002eaa",
  2700 => x"00001c9b",
  2701 => x"00000002",
  2702 => x"00002ec8",
  2703 => x"00001c9b",
  2704 => x"00000002",
  2705 => x"00002ee6",
  2706 => x"00001c9b",
  2707 => x"00000002",
  2708 => x"00002f04",
  2709 => x"00001c9b",
  2710 => x"00000002",
  2711 => x"00002f22",
  2712 => x"00001c9b",
  2713 => x"00000002",
  2714 => x"00002f40",
  2715 => x"00001c9b",
  2716 => x"00000002",
  2717 => x"00002f5e",
  2718 => x"00001c9b",
  2719 => x"00000002",
  2720 => x"00002f7c",
  2721 => x"00001c9b",
  2722 => x"00000002",
  2723 => x"00002f9a",
  2724 => x"00001c9b",
  2725 => x"00000002",
  2726 => x"00002fb8",
  2727 => x"00001c9b",
  2728 => x"00000002",
  2729 => x"00002fd6",
  2730 => x"00001c9b",
  2731 => x"00000002",
  2732 => x"00002ff4",
  2733 => x"00001c9b",
  2734 => x"00000004",
  2735 => x"000025e4",
  2736 => x"00000000",
  2737 => x"00000000",
  2738 => x"00000000",
  2739 => x"00001e4d",
  2740 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

