-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d5",
     9 => x"fc080b0b",
    10 => x"80d68008",
    11 => x"0b0b80d6",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d6840c0b",
    16 => x"0b80d680",
    17 => x"0c0b0b80",
    18 => x"d5fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbf98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d5fc70",
    57 => x"80e0bc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518add",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d6",
    65 => x"8c0c9f0b",
    66 => x"80d6900c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d69008ff",
    70 => x"0580d690",
    71 => x"0c80d690",
    72 => x"088025e8",
    73 => x"3880d68c",
    74 => x"08ff0580",
    75 => x"d68c0c80",
    76 => x"d68c0880",
    77 => x"25d03880",
    78 => x"0b80d690",
    79 => x"0c800b80",
    80 => x"d68c0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d68c08",
   100 => x"25913882",
   101 => x"c82d80d6",
   102 => x"8c08ff05",
   103 => x"80d68c0c",
   104 => x"838a0480",
   105 => x"d68c0880",
   106 => x"d6900853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d68c08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d6900881",
   116 => x"0580d690",
   117 => x"0c80d690",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d690",
   121 => x"0c80d68c",
   122 => x"08810580",
   123 => x"d68c0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d6",
   128 => x"90088105",
   129 => x"80d6900c",
   130 => x"80d69008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d690",
   134 => x"0c80d68c",
   135 => x"08810580",
   136 => x"d68c0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d6940cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d6940c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d6",
   177 => x"94088407",
   178 => x"80d6940c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5483f474",
   182 => x"258f3883",
   183 => x"0b0b0b80",
   184 => x"cc940c82",
   185 => x"985385f3",
   186 => x"04810b0b",
   187 => x"0b80cc94",
   188 => x"0ca8530b",
   189 => x"0b80cc94",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0c747431",
   193 => x"ffb005ff",
   194 => x"1271712c",
   195 => x"ff941970",
   196 => x"9f2a1170",
   197 => x"812c80d6",
   198 => x"94085255",
   199 => x"51525652",
   200 => x"53517680",
   201 => x"2e853870",
   202 => x"81075170",
   203 => x"f6940c72",
   204 => x"098105f6",
   205 => x"800c7109",
   206 => x"8105f684",
   207 => x"0c029405",
   208 => x"0d040402",
   209 => x"fc050d80",
   210 => x"d2a05195",
   211 => x"cb2d0284",
   212 => x"050d0402",
   213 => x"fc050d80",
   214 => x"cc985195",
   215 => x"cb2d0284",
   216 => x"050d0402",
   217 => x"fc050d80",
   218 => x"d0f85195",
   219 => x"cb2d0284",
   220 => x"050d0402",
   221 => x"fc050d81",
   222 => x"808051c0",
   223 => x"115170fb",
   224 => x"38028405",
   225 => x"0d047181",
   226 => x"2e098106",
   227 => x"893881c3",
   228 => x"0bec0c87",
   229 => x"9a04830b",
   230 => x"ec0c86f3",
   231 => x"2d820bec",
   232 => x"0c049388",
   233 => x"2d80d5fc",
   234 => x"0880d0e8",
   235 => x"0c93882d",
   236 => x"80d5fc08",
   237 => x"80d0940c",
   238 => x"93882d80",
   239 => x"d5fc0880",
   240 => x"d3b80c93",
   241 => x"882d80d5",
   242 => x"fc0880d2",
   243 => x"900c9388",
   244 => x"2d80d5fc",
   245 => x"0880cdbc",
   246 => x"0c0402fc",
   247 => x"050d84bf",
   248 => x"5186f32d",
   249 => x"ff115170",
   250 => x"8025f638",
   251 => x"0284050d",
   252 => x"0402f405",
   253 => x"0d745372",
   254 => x"70810554",
   255 => x"80f52d52",
   256 => x"71802e89",
   257 => x"38715183",
   258 => x"842d87f7",
   259 => x"04810b80",
   260 => x"d5fc0c02",
   261 => x"8c050d04",
   262 => x"02dc050d",
   263 => x"800b80ce",
   264 => x"8c085459",
   265 => x"72822e89",
   266 => x"3872832e",
   267 => x"963888d5",
   268 => x"0480d6a4",
   269 => x"08bffaff",
   270 => x"06828007",
   271 => x"80d6a40c",
   272 => x"88e40480",
   273 => x"d6a408bf",
   274 => x"ffff0687",
   275 => x"800780d6",
   276 => x"a40c88e4",
   277 => x"0480d6a4",
   278 => x"08bff9ff",
   279 => x"06818007",
   280 => x"80d6a40c",
   281 => x"80d6a408",
   282 => x"fc0c8184",
   283 => x"0bec0c7a",
   284 => x"5280d698",
   285 => x"51b4c12d",
   286 => x"80d5fc08",
   287 => x"802e819d",
   288 => x"3880d69c",
   289 => x"08548056",
   290 => x"73852e09",
   291 => x"81068a38",
   292 => x"840bec0c",
   293 => x"81538aa5",
   294 => x"0473f80c",
   295 => x"81a40bec",
   296 => x"0c87da2d",
   297 => x"75ff1557",
   298 => x"5875802e",
   299 => x"8b388118",
   300 => x"76812a57",
   301 => x"5889a904",
   302 => x"f7185881",
   303 => x"59807425",
   304 => x"80d738a4",
   305 => x"0bec0c77",
   306 => x"52755184",
   307 => x"a82d80d6",
   308 => x"f45280d6",
   309 => x"9851b7b4",
   310 => x"2d80d5fc",
   311 => x"08802ea0",
   312 => x"3880d6f4",
   313 => x"5783fc55",
   314 => x"76708405",
   315 => x"5808e80c",
   316 => x"fc155574",
   317 => x"8025f138",
   318 => x"81a40bec",
   319 => x"0c8a8804",
   320 => x"80d5fc08",
   321 => x"59848054",
   322 => x"80d69851",
   323 => x"b7842dfc",
   324 => x"80148117",
   325 => x"575489bd",
   326 => x"04840bec",
   327 => x"0c80d69c",
   328 => x"08f80c78",
   329 => x"537280d5",
   330 => x"fc0c02a4",
   331 => x"050d0402",
   332 => x"f8050d73",
   333 => x"5188982d",
   334 => x"80d5fc08",
   335 => x"5280d5fc",
   336 => x"08802e88",
   337 => x"3880d0a4",
   338 => x"518ad004",
   339 => x"80d08051",
   340 => x"95cb2d71",
   341 => x"80d5fc0c",
   342 => x"0288050d",
   343 => x"0402f005",
   344 => x"0d800b80",
   345 => x"d6a40c81",
   346 => x"5187862d",
   347 => x"80518786",
   348 => x"2d840bec",
   349 => x"0c92d82d",
   350 => x"8f832d81",
   351 => x"f92d8352",
   352 => x"92bb2d81",
   353 => x"51858d2d",
   354 => x"ff125271",
   355 => x"8025f138",
   356 => x"80c40bec",
   357 => x"0c80c9e8",
   358 => x"5187f12d",
   359 => x"aaf92d80",
   360 => x"d5fc0880",
   361 => x"2e83c538",
   362 => x"81840bec",
   363 => x"0c80ca80",
   364 => x"5187f12d",
   365 => x"80d6a408",
   366 => x"bfffff06",
   367 => x"87800770",
   368 => x"80d6a40c",
   369 => x"fc0c80ca",
   370 => x"98518898",
   371 => x"2d80d5fc",
   372 => x"08802e80",
   373 => x"cc3880ca",
   374 => x"a4518898",
   375 => x"2d80d5fc",
   376 => x"08802ebd",
   377 => x"3880cab0",
   378 => x"5188982d",
   379 => x"80d5fc08",
   380 => x"5280d5fc",
   381 => x"08973880",
   382 => x"cabc5187",
   383 => x"f12d80ca",
   384 => x"d4518898",
   385 => x"2d715187",
   386 => x"862d8ca8",
   387 => x"0480cad4",
   388 => x"5188982d",
   389 => x"80518786",
   390 => x"2d805185",
   391 => x"8d2d8ca8",
   392 => x"0480cabc",
   393 => x"5187f12d",
   394 => x"840bec0c",
   395 => x"8aaf51bf",
   396 => x"902d80d6",
   397 => x"a40880d4",
   398 => x"900c80d6",
   399 => x"a408fc0c",
   400 => x"80d6d408",
   401 => x"882a7081",
   402 => x"06515271",
   403 => x"802e8c38",
   404 => x"80cf880b",
   405 => x"80d6a80c",
   406 => x"8ce30480",
   407 => x"ce900b80",
   408 => x"d6a80c80",
   409 => x"d6a80851",
   410 => x"95cb2d80",
   411 => x"5187a22d",
   412 => x"830b80d6",
   413 => x"e80c9391",
   414 => x"2d805185",
   415 => x"8d2d93a5",
   416 => x"2d8f8f2d",
   417 => x"95de2d80",
   418 => x"ccb80b80",
   419 => x"f52d80cc",
   420 => x"c40b80f5",
   421 => x"2d718a2b",
   422 => x"718b2b07",
   423 => x"80ccdc0b",
   424 => x"80f52d70",
   425 => x"8d2b7207",
   426 => x"80ccf40b",
   427 => x"80f52d70",
   428 => x"8e2b7207",
   429 => x"80cda40b",
   430 => x"80f52d70",
   431 => x"912b7207",
   432 => x"7080d6a4",
   433 => x"0c80d490",
   434 => x"08708106",
   435 => x"54525354",
   436 => x"52545253",
   437 => x"54555371",
   438 => x"802e8838",
   439 => x"73810780",
   440 => x"d6a40c72",
   441 => x"812a7081",
   442 => x"06515271",
   443 => x"802e8b38",
   444 => x"80d6a408",
   445 => x"820780d6",
   446 => x"a40c7282",
   447 => x"2a708106",
   448 => x"51527180",
   449 => x"2e8b3880",
   450 => x"d6a40884",
   451 => x"0780d6a4",
   452 => x"0c72832a",
   453 => x"70810651",
   454 => x"5271802e",
   455 => x"8b3880d6",
   456 => x"a4088807",
   457 => x"80d6a40c",
   458 => x"72842a70",
   459 => x"81065152",
   460 => x"71802e8b",
   461 => x"3880d6a4",
   462 => x"08900780",
   463 => x"d6a40c72",
   464 => x"852a7081",
   465 => x"06515271",
   466 => x"802e8b38",
   467 => x"80d6a408",
   468 => x"a00780d6",
   469 => x"a40c80d6",
   470 => x"a408fc0c",
   471 => x"865280d5",
   472 => x"fc088338",
   473 => x"845271ec",
   474 => x"0c8d8104",
   475 => x"800b80d5",
   476 => x"fc0c0290",
   477 => x"050d0471",
   478 => x"980c04ff",
   479 => x"b00880d5",
   480 => x"fc0c0481",
   481 => x"0bffb00c",
   482 => x"04800bff",
   483 => x"b00c0402",
   484 => x"f4050d90",
   485 => x"9d0480d5",
   486 => x"fc0881f0",
   487 => x"2e098106",
   488 => x"8a38810b",
   489 => x"80d4880c",
   490 => x"909d0480",
   491 => x"d5fc0881",
   492 => x"e02e0981",
   493 => x"068a3881",
   494 => x"0b80d48c",
   495 => x"0c909d04",
   496 => x"80d5fc08",
   497 => x"5280d48c",
   498 => x"08802e89",
   499 => x"3880d5fc",
   500 => x"08818005",
   501 => x"5271842c",
   502 => x"728f0653",
   503 => x"5380d488",
   504 => x"08802e9a",
   505 => x"38728429",
   506 => x"80d3c805",
   507 => x"72138171",
   508 => x"2b700973",
   509 => x"0806730c",
   510 => x"51535390",
   511 => x"91047284",
   512 => x"2980d3c8",
   513 => x"05721383",
   514 => x"712b7208",
   515 => x"07720c53",
   516 => x"53800b80",
   517 => x"d48c0c80",
   518 => x"0b80d488",
   519 => x"0c80d6ac",
   520 => x"5191a42d",
   521 => x"80d5fc08",
   522 => x"ff24feea",
   523 => x"38800b80",
   524 => x"d5fc0c02",
   525 => x"8c050d04",
   526 => x"02f8050d",
   527 => x"80d3c852",
   528 => x"8f518072",
   529 => x"70840554",
   530 => x"0cff1151",
   531 => x"708025f2",
   532 => x"38028805",
   533 => x"0d0402f0",
   534 => x"050d7551",
   535 => x"8f892d70",
   536 => x"822cfc06",
   537 => x"80d3c811",
   538 => x"72109e06",
   539 => x"71087072",
   540 => x"2a708306",
   541 => x"82742b70",
   542 => x"09740676",
   543 => x"0c545156",
   544 => x"57535153",
   545 => x"8f832d71",
   546 => x"80d5fc0c",
   547 => x"0290050d",
   548 => x"0402fc05",
   549 => x"0d725180",
   550 => x"710c800b",
   551 => x"84120c02",
   552 => x"84050d04",
   553 => x"02f0050d",
   554 => x"75700884",
   555 => x"12085353",
   556 => x"53ff5471",
   557 => x"712ea838",
   558 => x"8f892d84",
   559 => x"13087084",
   560 => x"29148811",
   561 => x"70087081",
   562 => x"ff068418",
   563 => x"08811187",
   564 => x"06841a0c",
   565 => x"53515551",
   566 => x"51518f83",
   567 => x"2d715473",
   568 => x"80d5fc0c",
   569 => x"0290050d",
   570 => x"0402f405",
   571 => x"0d8f892d",
   572 => x"e008708b",
   573 => x"2a708106",
   574 => x"51525370",
   575 => x"802ea138",
   576 => x"80d6ac08",
   577 => x"70842980",
   578 => x"d6b40574",
   579 => x"81ff0671",
   580 => x"0c515180",
   581 => x"d6ac0881",
   582 => x"11870680",
   583 => x"d6ac0c51",
   584 => x"728c2c83",
   585 => x"ff0680d6",
   586 => x"d40c800b",
   587 => x"80d6d80c",
   588 => x"8efb2d8f",
   589 => x"832d028c",
   590 => x"050d0402",
   591 => x"fc050d8f",
   592 => x"892d810b",
   593 => x"80d6d80c",
   594 => x"8f832d80",
   595 => x"d6d80851",
   596 => x"70f93802",
   597 => x"84050d04",
   598 => x"02fc050d",
   599 => x"80d6ac51",
   600 => x"91912d90",
   601 => x"b82d91e9",
   602 => x"518ef72d",
   603 => x"0284050d",
   604 => x"0402fc05",
   605 => x"0d8fcf51",
   606 => x"86f32dff",
   607 => x"11517080",
   608 => x"25f63802",
   609 => x"84050d04",
   610 => x"80d6e008",
   611 => x"80d5fc0c",
   612 => x"0402fc05",
   613 => x"0d810b80",
   614 => x"d4bc0c81",
   615 => x"51858d2d",
   616 => x"0284050d",
   617 => x"0402fc05",
   618 => x"0d93af04",
   619 => x"8f8f2d80",
   620 => x"f65190d6",
   621 => x"2d80d5fc",
   622 => x"08f23880",
   623 => x"da5190d6",
   624 => x"2d80d5fc",
   625 => x"08e63880",
   626 => x"d4b80851",
   627 => x"90d62d80",
   628 => x"d5fc08d8",
   629 => x"38835190",
   630 => x"d62d80d5",
   631 => x"fc08cd38",
   632 => x"80d5fc08",
   633 => x"80d4bc0c",
   634 => x"80d5fc08",
   635 => x"51858d2d",
   636 => x"0284050d",
   637 => x"0402ec05",
   638 => x"0d765480",
   639 => x"52870b88",
   640 => x"1580f52d",
   641 => x"56537472",
   642 => x"248338a0",
   643 => x"53725183",
   644 => x"842d8112",
   645 => x"8b1580f5",
   646 => x"2d545272",
   647 => x"7225de38",
   648 => x"0294050d",
   649 => x"0402f005",
   650 => x"0d80d6e0",
   651 => x"085481f9",
   652 => x"2d800b80",
   653 => x"d6e40c73",
   654 => x"08802e81",
   655 => x"8938820b",
   656 => x"80d6900c",
   657 => x"80d6e408",
   658 => x"8f0680d6",
   659 => x"8c0c7308",
   660 => x"5271832e",
   661 => x"96387183",
   662 => x"26893871",
   663 => x"812eb038",
   664 => x"95af0471",
   665 => x"852ea038",
   666 => x"95af0488",
   667 => x"1480f52d",
   668 => x"84150880",
   669 => x"cae05354",
   670 => x"5287f12d",
   671 => x"71842913",
   672 => x"70085252",
   673 => x"95b30473",
   674 => x"5193f52d",
   675 => x"95af0480",
   676 => x"d4900888",
   677 => x"15082c70",
   678 => x"81065152",
   679 => x"71802e88",
   680 => x"3880cae4",
   681 => x"5195ac04",
   682 => x"80cae851",
   683 => x"87f12d84",
   684 => x"14085187",
   685 => x"f12d80d6",
   686 => x"e4088105",
   687 => x"80d6e40c",
   688 => x"8c145494",
   689 => x"b7040290",
   690 => x"050d0471",
   691 => x"80d6e00c",
   692 => x"94a52d80",
   693 => x"d6e408ff",
   694 => x"0580d6e8",
   695 => x"0c0402e8",
   696 => x"050d80d6",
   697 => x"e00880d6",
   698 => x"ec085755",
   699 => x"80f65190",
   700 => x"d62d80d5",
   701 => x"fc08812a",
   702 => x"70810651",
   703 => x"52719c38",
   704 => x"835190d6",
   705 => x"2d80d5fc",
   706 => x"08812a70",
   707 => x"81065152",
   708 => x"71802ead",
   709 => x"38969b04",
   710 => x"8f8f2d80",
   711 => x"f65190d6",
   712 => x"2d80d5fc",
   713 => x"08f23883",
   714 => x"5190d62d",
   715 => x"80d5fc08",
   716 => x"e73880d4",
   717 => x"bc088132",
   718 => x"7080d4bc",
   719 => x"0c51858d",
   720 => x"2d800b80",
   721 => x"d6dc0c8c",
   722 => x"5190d62d",
   723 => x"80d5fc08",
   724 => x"812a7081",
   725 => x"06515271",
   726 => x"802e80d1",
   727 => x"3880d494",
   728 => x"0880d4a8",
   729 => x"0880d494",
   730 => x"0c80d4a8",
   731 => x"0c80d498",
   732 => x"0880d4ac",
   733 => x"0880d498",
   734 => x"0c80d4ac",
   735 => x"0c80d49c",
   736 => x"0880d4b0",
   737 => x"0880d49c",
   738 => x"0c80d4b0",
   739 => x"0c80d4a0",
   740 => x"0880d4b4",
   741 => x"0880d4a0",
   742 => x"0c80d4b4",
   743 => x"0c80d4a4",
   744 => x"0880d4b8",
   745 => x"0880d4a4",
   746 => x"0c80d4b8",
   747 => x"0c80d6d4",
   748 => x"08a00652",
   749 => x"80722596",
   750 => x"3892f12d",
   751 => x"8f8f2d80",
   752 => x"d4bc0881",
   753 => x"327080d4",
   754 => x"bc0c5185",
   755 => x"8d2d80d4",
   756 => x"bc0882ef",
   757 => x"3880d4a8",
   758 => x"085190d6",
   759 => x"2d80d5fc",
   760 => x"08802e8b",
   761 => x"3880d6dc",
   762 => x"08810780",
   763 => x"d6dc0c80",
   764 => x"d4ac0851",
   765 => x"90d62d80",
   766 => x"d5fc0880",
   767 => x"2e8b3880",
   768 => x"d6dc0882",
   769 => x"0780d6dc",
   770 => x"0c80d4b0",
   771 => x"085190d6",
   772 => x"2d80d5fc",
   773 => x"08802e8b",
   774 => x"3880d6dc",
   775 => x"08840780",
   776 => x"d6dc0c80",
   777 => x"d4b40851",
   778 => x"90d62d80",
   779 => x"d5fc0880",
   780 => x"2e8b3880",
   781 => x"d6dc0888",
   782 => x"0780d6dc",
   783 => x"0c80d4b8",
   784 => x"085190d6",
   785 => x"2d80d5fc",
   786 => x"08802e8b",
   787 => x"3880d6dc",
   788 => x"08900780",
   789 => x"d6dc0c80",
   790 => x"d4940851",
   791 => x"90d62d80",
   792 => x"d5fc0880",
   793 => x"2e8c3880",
   794 => x"d6dc0882",
   795 => x"800780d6",
   796 => x"dc0c80d4",
   797 => x"98085190",
   798 => x"d62d80d5",
   799 => x"fc08802e",
   800 => x"8c3880d6",
   801 => x"dc088480",
   802 => x"0780d6dc",
   803 => x"0c80d49c",
   804 => x"085190d6",
   805 => x"2d80d5fc",
   806 => x"08802e8c",
   807 => x"3880d6dc",
   808 => x"08888007",
   809 => x"80d6dc0c",
   810 => x"80d4a008",
   811 => x"5190d62d",
   812 => x"80d5fc08",
   813 => x"802e8c38",
   814 => x"80d6dc08",
   815 => x"90800780",
   816 => x"d6dc0c80",
   817 => x"d4a40851",
   818 => x"90d62d80",
   819 => x"d5fc0880",
   820 => x"2e8c3880",
   821 => x"d6dc08a0",
   822 => x"800780d6",
   823 => x"dc0c9451",
   824 => x"90d62d80",
   825 => x"d5fc0852",
   826 => x"915190d6",
   827 => x"2d7180d5",
   828 => x"fc080652",
   829 => x"80e65190",
   830 => x"d62d7180",
   831 => x"d5fc0806",
   832 => x"5271802e",
   833 => x"8d3880d6",
   834 => x"dc088480",
   835 => x"800780d6",
   836 => x"dc0c80fe",
   837 => x"5190d62d",
   838 => x"80d5fc08",
   839 => x"52875190",
   840 => x"d62d7180",
   841 => x"d5fc0807",
   842 => x"5271802e",
   843 => x"8d3880d6",
   844 => x"dc088880",
   845 => x"800780d6",
   846 => x"dc0c80d6",
   847 => x"dc08ed0c",
   848 => x"a2ce0494",
   849 => x"5190d62d",
   850 => x"80d5fc08",
   851 => x"52915190",
   852 => x"d62d7180",
   853 => x"d5fc0806",
   854 => x"5280e651",
   855 => x"90d62d71",
   856 => x"80d5fc08",
   857 => x"06527180",
   858 => x"2e8d3880",
   859 => x"d6dc0884",
   860 => x"80800780",
   861 => x"d6dc0c80",
   862 => x"fe5190d6",
   863 => x"2d80d5fc",
   864 => x"08528751",
   865 => x"90d62d71",
   866 => x"80d5fc08",
   867 => x"07527180",
   868 => x"2e8d3880",
   869 => x"d6dc0888",
   870 => x"80800780",
   871 => x"d6dc0c80",
   872 => x"d6dc08ed",
   873 => x"0c81f551",
   874 => x"90d62d80",
   875 => x"d5fc0881",
   876 => x"2a708106",
   877 => x"515271a4",
   878 => x"3880d4a8",
   879 => x"085190d6",
   880 => x"2d80d5fc",
   881 => x"08812a70",
   882 => x"81065152",
   883 => x"718e3880",
   884 => x"d6d40881",
   885 => x"06528072",
   886 => x"2580c238",
   887 => x"80d6d408",
   888 => x"81065280",
   889 => x"72258438",
   890 => x"92f12d80",
   891 => x"d6e80852",
   892 => x"71802e8a",
   893 => x"38ff1280",
   894 => x"d6e80c9c",
   895 => x"9d0480d6",
   896 => x"e4081080",
   897 => x"d6e40805",
   898 => x"70842916",
   899 => x"51528812",
   900 => x"08802e89",
   901 => x"38ff5188",
   902 => x"12085271",
   903 => x"2d81f251",
   904 => x"90d62d80",
   905 => x"d5fc0881",
   906 => x"2a708106",
   907 => x"515271a4",
   908 => x"3880d4ac",
   909 => x"085190d6",
   910 => x"2d80d5fc",
   911 => x"08812a70",
   912 => x"81065152",
   913 => x"718e3880",
   914 => x"d6d40882",
   915 => x"06528072",
   916 => x"2580c338",
   917 => x"80d6d408",
   918 => x"82065280",
   919 => x"72258438",
   920 => x"92f12d80",
   921 => x"d6e408ff",
   922 => x"1180d6e8",
   923 => x"08565353",
   924 => x"7372258a",
   925 => x"38811480",
   926 => x"d6e80c9d",
   927 => x"96047210",
   928 => x"13708429",
   929 => x"16515288",
   930 => x"1208802e",
   931 => x"8938fe51",
   932 => x"88120852",
   933 => x"712d81fd",
   934 => x"5190d62d",
   935 => x"80d5fc08",
   936 => x"812a7081",
   937 => x"06515271",
   938 => x"a43880d4",
   939 => x"b0085190",
   940 => x"d62d80d5",
   941 => x"fc08812a",
   942 => x"70810651",
   943 => x"52718e38",
   944 => x"80d6d408",
   945 => x"84065280",
   946 => x"722580c0",
   947 => x"3880d6d4",
   948 => x"08840652",
   949 => x"80722584",
   950 => x"3892f12d",
   951 => x"80d6e808",
   952 => x"802e8a38",
   953 => x"800b80d6",
   954 => x"e80c9e8c",
   955 => x"0480d6e4",
   956 => x"081080d6",
   957 => x"e4080570",
   958 => x"84291651",
   959 => x"52881208",
   960 => x"802e8938",
   961 => x"fd518812",
   962 => x"0852712d",
   963 => x"81fa5190",
   964 => x"d62d80d5",
   965 => x"fc08812a",
   966 => x"70810651",
   967 => x"5271a438",
   968 => x"80d4b408",
   969 => x"5190d62d",
   970 => x"80d5fc08",
   971 => x"812a7081",
   972 => x"06515271",
   973 => x"8e3880d6",
   974 => x"d4088806",
   975 => x"52807225",
   976 => x"80c03880",
   977 => x"d6d40888",
   978 => x"06528072",
   979 => x"25843892",
   980 => x"f12d80d6",
   981 => x"e408ff11",
   982 => x"545280d6",
   983 => x"e8087325",
   984 => x"89387280",
   985 => x"d6e80c9f",
   986 => x"82047110",
   987 => x"12708429",
   988 => x"16515288",
   989 => x"1208802e",
   990 => x"8938fc51",
   991 => x"88120852",
   992 => x"712d80d6",
   993 => x"e8087053",
   994 => x"5473802e",
   995 => x"8a388c15",
   996 => x"ff155555",
   997 => x"9f890482",
   998 => x"0b80d690",
   999 => x"0c718f06",
  1000 => x"80d68c0c",
  1001 => x"81eb5190",
  1002 => x"d62d80d5",
  1003 => x"fc08812a",
  1004 => x"70810651",
  1005 => x"5271802e",
  1006 => x"ad387408",
  1007 => x"852e0981",
  1008 => x"06a43888",
  1009 => x"1580f52d",
  1010 => x"ff055271",
  1011 => x"881681b7",
  1012 => x"2d71982b",
  1013 => x"52718025",
  1014 => x"8838800b",
  1015 => x"881681b7",
  1016 => x"2d745193",
  1017 => x"f52d81f4",
  1018 => x"5190d62d",
  1019 => x"80d5fc08",
  1020 => x"812a7081",
  1021 => x"06515271",
  1022 => x"802eb338",
  1023 => x"7408852e",
  1024 => x"098106aa",
  1025 => x"38881580",
  1026 => x"f52d8105",
  1027 => x"52718816",
  1028 => x"81b72d71",
  1029 => x"81ff068b",
  1030 => x"1680f52d",
  1031 => x"54527272",
  1032 => x"27873872",
  1033 => x"881681b7",
  1034 => x"2d745193",
  1035 => x"f52d80da",
  1036 => x"5190d62d",
  1037 => x"80d5fc08",
  1038 => x"812a7081",
  1039 => x"06515271",
  1040 => x"8e3880d6",
  1041 => x"d4089006",
  1042 => x"52807225",
  1043 => x"81bc3880",
  1044 => x"d6e00880",
  1045 => x"d6d40890",
  1046 => x"06535380",
  1047 => x"72258438",
  1048 => x"92f12d80",
  1049 => x"d6e80854",
  1050 => x"73802e8a",
  1051 => x"388c13ff",
  1052 => x"155553a0",
  1053 => x"e8047208",
  1054 => x"5271822e",
  1055 => x"a6387182",
  1056 => x"26893871",
  1057 => x"812eaa38",
  1058 => x"a28a0471",
  1059 => x"832eb438",
  1060 => x"71842e09",
  1061 => x"810680f2",
  1062 => x"38881308",
  1063 => x"5195cb2d",
  1064 => x"a28a0480",
  1065 => x"d6e80851",
  1066 => x"88130852",
  1067 => x"712da28a",
  1068 => x"04810b88",
  1069 => x"14082b80",
  1070 => x"d4900832",
  1071 => x"80d4900c",
  1072 => x"a1de0488",
  1073 => x"1380f52d",
  1074 => x"81058b14",
  1075 => x"80f52d53",
  1076 => x"54717424",
  1077 => x"83388054",
  1078 => x"73881481",
  1079 => x"b72d94a5",
  1080 => x"2da28a04",
  1081 => x"7508802e",
  1082 => x"a4387508",
  1083 => x"5190d62d",
  1084 => x"80d5fc08",
  1085 => x"81065271",
  1086 => x"802e8c38",
  1087 => x"80d6e808",
  1088 => x"51841608",
  1089 => x"52712d88",
  1090 => x"165675d8",
  1091 => x"38805480",
  1092 => x"0b80d690",
  1093 => x"0c738f06",
  1094 => x"80d68c0c",
  1095 => x"a0527380",
  1096 => x"d6e8082e",
  1097 => x"09810699",
  1098 => x"3880d6e4",
  1099 => x"08ff0574",
  1100 => x"32700981",
  1101 => x"05707207",
  1102 => x"9f2a9171",
  1103 => x"31515153",
  1104 => x"53715183",
  1105 => x"842d8114",
  1106 => x"548e7425",
  1107 => x"c23880d4",
  1108 => x"bc0880d5",
  1109 => x"fc0c0298",
  1110 => x"050d0402",
  1111 => x"f4050dd4",
  1112 => x"5281ff72",
  1113 => x"0c710853",
  1114 => x"81ff720c",
  1115 => x"72882b83",
  1116 => x"fe800672",
  1117 => x"087081ff",
  1118 => x"06515253",
  1119 => x"81ff720c",
  1120 => x"72710788",
  1121 => x"2b720870",
  1122 => x"81ff0651",
  1123 => x"525381ff",
  1124 => x"720c7271",
  1125 => x"07882b72",
  1126 => x"087081ff",
  1127 => x"06720780",
  1128 => x"d5fc0c52",
  1129 => x"53028c05",
  1130 => x"0d0402f4",
  1131 => x"050d7476",
  1132 => x"7181ff06",
  1133 => x"d40c5353",
  1134 => x"80d6f008",
  1135 => x"85387189",
  1136 => x"2b527198",
  1137 => x"2ad40c71",
  1138 => x"902a7081",
  1139 => x"ff06d40c",
  1140 => x"5171882a",
  1141 => x"7081ff06",
  1142 => x"d40c5171",
  1143 => x"81ff06d4",
  1144 => x"0c72902a",
  1145 => x"7081ff06",
  1146 => x"d40c51d4",
  1147 => x"087081ff",
  1148 => x"06515182",
  1149 => x"b8bf5270",
  1150 => x"81ff2e09",
  1151 => x"81069438",
  1152 => x"81ff0bd4",
  1153 => x"0cd40870",
  1154 => x"81ff06ff",
  1155 => x"14545151",
  1156 => x"71e53870",
  1157 => x"80d5fc0c",
  1158 => x"028c050d",
  1159 => x"0402fc05",
  1160 => x"0d81c751",
  1161 => x"81ff0bd4",
  1162 => x"0cff1151",
  1163 => x"708025f4",
  1164 => x"38028405",
  1165 => x"0d0402f4",
  1166 => x"050d81ff",
  1167 => x"0bd40c93",
  1168 => x"53805287",
  1169 => x"fc80c151",
  1170 => x"a3aa2d80",
  1171 => x"d5fc088b",
  1172 => x"3881ff0b",
  1173 => x"d40c8153",
  1174 => x"a4e404a4",
  1175 => x"9d2dff13",
  1176 => x"5372de38",
  1177 => x"7280d5fc",
  1178 => x"0c028c05",
  1179 => x"0d0402ec",
  1180 => x"050d810b",
  1181 => x"80d6f00c",
  1182 => x"8454d008",
  1183 => x"708f2a70",
  1184 => x"81065151",
  1185 => x"5372f338",
  1186 => x"72d00ca4",
  1187 => x"9d2d80ca",
  1188 => x"ec5187f1",
  1189 => x"2dd00870",
  1190 => x"8f2a7081",
  1191 => x"06515153",
  1192 => x"72f33881",
  1193 => x"0bd00cb1",
  1194 => x"53805284",
  1195 => x"d480c051",
  1196 => x"a3aa2d80",
  1197 => x"d5fc0881",
  1198 => x"2e933872",
  1199 => x"822ebf38",
  1200 => x"ff135372",
  1201 => x"e438ff14",
  1202 => x"5473ffae",
  1203 => x"38a49d2d",
  1204 => x"83aa5284",
  1205 => x"9c80c851",
  1206 => x"a3aa2d80",
  1207 => x"d5fc0881",
  1208 => x"2e098106",
  1209 => x"9338a2db",
  1210 => x"2d80d5fc",
  1211 => x"0883ffff",
  1212 => x"06537283",
  1213 => x"aa2e9f38",
  1214 => x"a4b62da6",
  1215 => x"910480ca",
  1216 => x"f85187f1",
  1217 => x"2d8053a7",
  1218 => x"e60480cb",
  1219 => x"905187f1",
  1220 => x"2d8054a7",
  1221 => x"b70481ff",
  1222 => x"0bd40cb1",
  1223 => x"54a49d2d",
  1224 => x"8fcf5380",
  1225 => x"5287fc80",
  1226 => x"f751a3aa",
  1227 => x"2d80d5fc",
  1228 => x"085580d5",
  1229 => x"fc08812e",
  1230 => x"0981069c",
  1231 => x"3881ff0b",
  1232 => x"d40c820a",
  1233 => x"52849c80",
  1234 => x"e951a3aa",
  1235 => x"2d80d5fc",
  1236 => x"08802e8d",
  1237 => x"38a49d2d",
  1238 => x"ff135372",
  1239 => x"c638a7aa",
  1240 => x"0481ff0b",
  1241 => x"d40c80d5",
  1242 => x"fc085287",
  1243 => x"fc80fa51",
  1244 => x"a3aa2d80",
  1245 => x"d5fc08b2",
  1246 => x"3881ff0b",
  1247 => x"d40cd408",
  1248 => x"5381ff0b",
  1249 => x"d40c81ff",
  1250 => x"0bd40c81",
  1251 => x"ff0bd40c",
  1252 => x"81ff0bd4",
  1253 => x"0c72862a",
  1254 => x"70810676",
  1255 => x"56515372",
  1256 => x"963880d5",
  1257 => x"fc0854a7",
  1258 => x"b7047382",
  1259 => x"2efedb38",
  1260 => x"ff145473",
  1261 => x"fee73873",
  1262 => x"80d6f00c",
  1263 => x"738b3881",
  1264 => x"5287fc80",
  1265 => x"d051a3aa",
  1266 => x"2d81ff0b",
  1267 => x"d40cd008",
  1268 => x"708f2a70",
  1269 => x"81065151",
  1270 => x"5372f338",
  1271 => x"72d00c81",
  1272 => x"ff0bd40c",
  1273 => x"81537280",
  1274 => x"d5fc0c02",
  1275 => x"94050d04",
  1276 => x"02e8050d",
  1277 => x"78558056",
  1278 => x"81ff0bd4",
  1279 => x"0cd00870",
  1280 => x"8f2a7081",
  1281 => x"06515153",
  1282 => x"72f33882",
  1283 => x"810bd00c",
  1284 => x"81ff0bd4",
  1285 => x"0c775287",
  1286 => x"fc80d151",
  1287 => x"a3aa2d80",
  1288 => x"dbc6df54",
  1289 => x"80d5fc08",
  1290 => x"802e8b38",
  1291 => x"80cbb051",
  1292 => x"87f12da9",
  1293 => x"8a0481ff",
  1294 => x"0bd40cd4",
  1295 => x"087081ff",
  1296 => x"06515372",
  1297 => x"81fe2e09",
  1298 => x"81069e38",
  1299 => x"80ff53a2",
  1300 => x"db2d80d5",
  1301 => x"fc087570",
  1302 => x"8405570c",
  1303 => x"ff135372",
  1304 => x"8025ec38",
  1305 => x"8156a8ef",
  1306 => x"04ff1454",
  1307 => x"73c83881",
  1308 => x"ff0bd40c",
  1309 => x"81ff0bd4",
  1310 => x"0cd00870",
  1311 => x"8f2a7081",
  1312 => x"06515153",
  1313 => x"72f33872",
  1314 => x"d00c7580",
  1315 => x"d5fc0c02",
  1316 => x"98050d04",
  1317 => x"02e8050d",
  1318 => x"77797b58",
  1319 => x"55558053",
  1320 => x"727625a3",
  1321 => x"38747081",
  1322 => x"055680f5",
  1323 => x"2d747081",
  1324 => x"055680f5",
  1325 => x"2d525271",
  1326 => x"712e8638",
  1327 => x"8151a9c9",
  1328 => x"04811353",
  1329 => x"a9a00480",
  1330 => x"517080d5",
  1331 => x"fc0c0298",
  1332 => x"050d0402",
  1333 => x"ec050d76",
  1334 => x"5574802e",
  1335 => x"80c2389a",
  1336 => x"1580e02d",
  1337 => x"51b88e2d",
  1338 => x"80d5fc08",
  1339 => x"80d5fc08",
  1340 => x"80dda40c",
  1341 => x"80d5fc08",
  1342 => x"545480dd",
  1343 => x"8008802e",
  1344 => x"9a389415",
  1345 => x"80e02d51",
  1346 => x"b88e2d80",
  1347 => x"d5fc0890",
  1348 => x"2b83fff0",
  1349 => x"0a067075",
  1350 => x"07515372",
  1351 => x"80dda40c",
  1352 => x"80dda408",
  1353 => x"5372802e",
  1354 => x"9d3880dc",
  1355 => x"f808fe14",
  1356 => x"712980dd",
  1357 => x"8c080580",
  1358 => x"dda80c70",
  1359 => x"842b80dd",
  1360 => x"840c54aa",
  1361 => x"f40480dd",
  1362 => x"900880dd",
  1363 => x"a40c80dd",
  1364 => x"940880dd",
  1365 => x"a80c80dd",
  1366 => x"8008802e",
  1367 => x"8b3880dc",
  1368 => x"f808842b",
  1369 => x"53aaef04",
  1370 => x"80dd9808",
  1371 => x"842b5372",
  1372 => x"80dd840c",
  1373 => x"0294050d",
  1374 => x"0402d805",
  1375 => x"0d800b80",
  1376 => x"dd800c84",
  1377 => x"54a4ee2d",
  1378 => x"80d5fc08",
  1379 => x"802e9738",
  1380 => x"80d6f452",
  1381 => x"8051a7f0",
  1382 => x"2d80d5fc",
  1383 => x"08802e86",
  1384 => x"38fe54ab",
  1385 => x"ae04ff14",
  1386 => x"54738024",
  1387 => x"d838738d",
  1388 => x"3880cbc0",
  1389 => x"5187f12d",
  1390 => x"7355b183",
  1391 => x"04805681",
  1392 => x"0b80ddac",
  1393 => x"0c885380",
  1394 => x"cbd45280",
  1395 => x"d7aa51a9",
  1396 => x"942d80d5",
  1397 => x"fc08762e",
  1398 => x"09810689",
  1399 => x"3880d5fc",
  1400 => x"0880ddac",
  1401 => x"0c885380",
  1402 => x"cbe05280",
  1403 => x"d7c651a9",
  1404 => x"942d80d5",
  1405 => x"fc088938",
  1406 => x"80d5fc08",
  1407 => x"80ddac0c",
  1408 => x"80ddac08",
  1409 => x"802e8181",
  1410 => x"3880daba",
  1411 => x"0b80f52d",
  1412 => x"80dabb0b",
  1413 => x"80f52d71",
  1414 => x"982b7190",
  1415 => x"2b0780da",
  1416 => x"bc0b80f5",
  1417 => x"2d70882b",
  1418 => x"720780da",
  1419 => x"bd0b80f5",
  1420 => x"2d710780",
  1421 => x"daf20b80",
  1422 => x"f52d80da",
  1423 => x"f30b80f5",
  1424 => x"2d71882b",
  1425 => x"07535f54",
  1426 => x"525a5657",
  1427 => x"557381ab",
  1428 => x"aa2e0981",
  1429 => x"068e3875",
  1430 => x"51b7dd2d",
  1431 => x"80d5fc08",
  1432 => x"56acf204",
  1433 => x"7382d4d5",
  1434 => x"2e883880",
  1435 => x"cbec51ad",
  1436 => x"be0480d6",
  1437 => x"f4527551",
  1438 => x"a7f02d80",
  1439 => x"d5fc0855",
  1440 => x"80d5fc08",
  1441 => x"802e83fb",
  1442 => x"38885380",
  1443 => x"cbe05280",
  1444 => x"d7c651a9",
  1445 => x"942d80d5",
  1446 => x"fc088a38",
  1447 => x"810b80dd",
  1448 => x"800cadc4",
  1449 => x"04885380",
  1450 => x"cbd45280",
  1451 => x"d7aa51a9",
  1452 => x"942d80d5",
  1453 => x"fc08802e",
  1454 => x"8b3880cc",
  1455 => x"805187f1",
  1456 => x"2daea304",
  1457 => x"80daf20b",
  1458 => x"80f52d54",
  1459 => x"7380d52e",
  1460 => x"09810680",
  1461 => x"ce3880da",
  1462 => x"f30b80f5",
  1463 => x"2d547381",
  1464 => x"aa2e0981",
  1465 => x"06bd3880",
  1466 => x"0b80d6f4",
  1467 => x"0b80f52d",
  1468 => x"56547481",
  1469 => x"e92e8338",
  1470 => x"81547481",
  1471 => x"eb2e8c38",
  1472 => x"80557375",
  1473 => x"2e098106",
  1474 => x"82f93880",
  1475 => x"d6ff0b80",
  1476 => x"f52d5574",
  1477 => x"8e3880d7",
  1478 => x"800b80f5",
  1479 => x"2d547382",
  1480 => x"2e863880",
  1481 => x"55b18304",
  1482 => x"80d7810b",
  1483 => x"80f52d70",
  1484 => x"80dcf80c",
  1485 => x"ff0580dc",
  1486 => x"fc0c80d7",
  1487 => x"820b80f5",
  1488 => x"2d80d783",
  1489 => x"0b80f52d",
  1490 => x"58760577",
  1491 => x"82802905",
  1492 => x"7080dd88",
  1493 => x"0c80d784",
  1494 => x"0b80f52d",
  1495 => x"7080dd9c",
  1496 => x"0c80dd80",
  1497 => x"08595758",
  1498 => x"76802e81",
  1499 => x"b7388853",
  1500 => x"80cbe052",
  1501 => x"80d7c651",
  1502 => x"a9942d80",
  1503 => x"d5fc0882",
  1504 => x"823880dc",
  1505 => x"f8087084",
  1506 => x"2b80dd84",
  1507 => x"0c7080dd",
  1508 => x"980c80d7",
  1509 => x"990b80f5",
  1510 => x"2d80d798",
  1511 => x"0b80f52d",
  1512 => x"71828029",
  1513 => x"0580d79a",
  1514 => x"0b80f52d",
  1515 => x"70848080",
  1516 => x"291280d7",
  1517 => x"9b0b80f5",
  1518 => x"2d708180",
  1519 => x"0a291270",
  1520 => x"80dda00c",
  1521 => x"80dd9c08",
  1522 => x"712980dd",
  1523 => x"88080570",
  1524 => x"80dd8c0c",
  1525 => x"80d7a10b",
  1526 => x"80f52d80",
  1527 => x"d7a00b80",
  1528 => x"f52d7182",
  1529 => x"80290580",
  1530 => x"d7a20b80",
  1531 => x"f52d7084",
  1532 => x"80802912",
  1533 => x"80d7a30b",
  1534 => x"80f52d70",
  1535 => x"982b81f0",
  1536 => x"0a067205",
  1537 => x"7080dd90",
  1538 => x"0cfe117e",
  1539 => x"29770580",
  1540 => x"dd940c52",
  1541 => x"59524354",
  1542 => x"5e515259",
  1543 => x"525d5759",
  1544 => x"57b0fc04",
  1545 => x"80d7860b",
  1546 => x"80f52d80",
  1547 => x"d7850b80",
  1548 => x"f52d7182",
  1549 => x"80290570",
  1550 => x"80dd840c",
  1551 => x"70a02983",
  1552 => x"ff057089",
  1553 => x"2a7080dd",
  1554 => x"980c80d7",
  1555 => x"8b0b80f5",
  1556 => x"2d80d78a",
  1557 => x"0b80f52d",
  1558 => x"71828029",
  1559 => x"057080dd",
  1560 => x"a00c7b71",
  1561 => x"291e7080",
  1562 => x"dd940c7d",
  1563 => x"80dd900c",
  1564 => x"730580dd",
  1565 => x"8c0c555e",
  1566 => x"51515555",
  1567 => x"8051a9d3",
  1568 => x"2d815574",
  1569 => x"80d5fc0c",
  1570 => x"02a8050d",
  1571 => x"0402ec05",
  1572 => x"0d767087",
  1573 => x"2c7180ff",
  1574 => x"06555654",
  1575 => x"80dd8008",
  1576 => x"8a387388",
  1577 => x"2c7481ff",
  1578 => x"06545580",
  1579 => x"d6f45280",
  1580 => x"dd880815",
  1581 => x"51a7f02d",
  1582 => x"80d5fc08",
  1583 => x"5480d5fc",
  1584 => x"08802eb8",
  1585 => x"3880dd80",
  1586 => x"08802e9a",
  1587 => x"38728429",
  1588 => x"80d6f405",
  1589 => x"70085253",
  1590 => x"b7dd2d80",
  1591 => x"d5fc08f0",
  1592 => x"0a0653b1",
  1593 => x"fa047210",
  1594 => x"80d6f405",
  1595 => x"7080e02d",
  1596 => x"5253b88e",
  1597 => x"2d80d5fc",
  1598 => x"08537254",
  1599 => x"7380d5fc",
  1600 => x"0c029405",
  1601 => x"0d0402e0",
  1602 => x"050d7970",
  1603 => x"842c80dd",
  1604 => x"a8080571",
  1605 => x"8f065255",
  1606 => x"53728a38",
  1607 => x"80d6f452",
  1608 => x"7351a7f0",
  1609 => x"2d72a029",
  1610 => x"80d6f405",
  1611 => x"54807480",
  1612 => x"f52d5653",
  1613 => x"74732e83",
  1614 => x"38815374",
  1615 => x"81e52e81",
  1616 => x"f4388170",
  1617 => x"74065458",
  1618 => x"72802e81",
  1619 => x"e8388b14",
  1620 => x"80f52d70",
  1621 => x"832a7906",
  1622 => x"5856769b",
  1623 => x"3880d4c0",
  1624 => x"08537289",
  1625 => x"387280da",
  1626 => x"f40b81b7",
  1627 => x"2d7680d4",
  1628 => x"c00c7353",
  1629 => x"b4b70475",
  1630 => x"8f2e0981",
  1631 => x"0681b638",
  1632 => x"749f068d",
  1633 => x"2980dae7",
  1634 => x"11515381",
  1635 => x"1480f52d",
  1636 => x"73708105",
  1637 => x"5581b72d",
  1638 => x"831480f5",
  1639 => x"2d737081",
  1640 => x"055581b7",
  1641 => x"2d851480",
  1642 => x"f52d7370",
  1643 => x"81055581",
  1644 => x"b72d8714",
  1645 => x"80f52d73",
  1646 => x"70810555",
  1647 => x"81b72d89",
  1648 => x"1480f52d",
  1649 => x"73708105",
  1650 => x"5581b72d",
  1651 => x"8e1480f5",
  1652 => x"2d737081",
  1653 => x"055581b7",
  1654 => x"2d901480",
  1655 => x"f52d7370",
  1656 => x"81055581",
  1657 => x"b72d9214",
  1658 => x"80f52d73",
  1659 => x"70810555",
  1660 => x"81b72d94",
  1661 => x"1480f52d",
  1662 => x"73708105",
  1663 => x"5581b72d",
  1664 => x"961480f5",
  1665 => x"2d737081",
  1666 => x"055581b7",
  1667 => x"2d981480",
  1668 => x"f52d7370",
  1669 => x"81055581",
  1670 => x"b72d9c14",
  1671 => x"80f52d73",
  1672 => x"70810555",
  1673 => x"81b72d9e",
  1674 => x"1480f52d",
  1675 => x"7381b72d",
  1676 => x"7780d4c0",
  1677 => x"0c805372",
  1678 => x"80d5fc0c",
  1679 => x"02a0050d",
  1680 => x"0402cc05",
  1681 => x"0d7e605e",
  1682 => x"5b800b80",
  1683 => x"dda40880",
  1684 => x"dda80859",
  1685 => x"5d568059",
  1686 => x"80dd8408",
  1687 => x"792e81de",
  1688 => x"38788f06",
  1689 => x"a0175754",
  1690 => x"73913880",
  1691 => x"d6f45276",
  1692 => x"51811757",
  1693 => x"a7f02d80",
  1694 => x"d6f45680",
  1695 => x"7680f52d",
  1696 => x"56547474",
  1697 => x"2e833881",
  1698 => x"547481e5",
  1699 => x"2e81a338",
  1700 => x"81707506",
  1701 => x"555a7380",
  1702 => x"2e819738",
  1703 => x"8b1680f5",
  1704 => x"2d709806",
  1705 => x"59547780",
  1706 => x"e3388b53",
  1707 => x"7c527551",
  1708 => x"a9942d80",
  1709 => x"d5fc0880",
  1710 => x"f9389c16",
  1711 => x"0851b7dd",
  1712 => x"2d80d5fc",
  1713 => x"08841c0c",
  1714 => x"9a1680e0",
  1715 => x"2d51b88e",
  1716 => x"2d80d5fc",
  1717 => x"0880d5fc",
  1718 => x"08881d0c",
  1719 => x"80d5fc08",
  1720 => x"555580dd",
  1721 => x"8008802e",
  1722 => x"99389416",
  1723 => x"80e02d51",
  1724 => x"b88e2d80",
  1725 => x"d5fc0890",
  1726 => x"2b83fff0",
  1727 => x"0a067016",
  1728 => x"51547388",
  1729 => x"1c0c777b",
  1730 => x"0cb6ad04",
  1731 => x"73842a70",
  1732 => x"81065154",
  1733 => x"73802e9a",
  1734 => x"388b537c",
  1735 => x"527551a9",
  1736 => x"942d80d5",
  1737 => x"fc088b38",
  1738 => x"7551a9d3",
  1739 => x"2d7954b6",
  1740 => x"fa048119",
  1741 => x"5980dd84",
  1742 => x"087926fe",
  1743 => x"a43880dd",
  1744 => x"8008802e",
  1745 => x"b3387b51",
  1746 => x"b18d2d80",
  1747 => x"d5fc0880",
  1748 => x"d5fc0880",
  1749 => x"fffffff8",
  1750 => x"06555c73",
  1751 => x"80ffffff",
  1752 => x"f82e9538",
  1753 => x"80d5fc08",
  1754 => x"fe0580dc",
  1755 => x"f8082980",
  1756 => x"dd8c0805",
  1757 => x"57b4d604",
  1758 => x"80547380",
  1759 => x"d5fc0c02",
  1760 => x"b4050d04",
  1761 => x"02f4050d",
  1762 => x"74700881",
  1763 => x"05710c70",
  1764 => x"0880dcfc",
  1765 => x"08065353",
  1766 => x"718f3888",
  1767 => x"130851b1",
  1768 => x"8d2d80d5",
  1769 => x"fc088814",
  1770 => x"0c810b80",
  1771 => x"d5fc0c02",
  1772 => x"8c050d04",
  1773 => x"02f0050d",
  1774 => x"75881108",
  1775 => x"fe0580dc",
  1776 => x"f8082980",
  1777 => x"dd8c0811",
  1778 => x"720880dc",
  1779 => x"fc080605",
  1780 => x"79555354",
  1781 => x"54a7f02d",
  1782 => x"0290050d",
  1783 => x"0402f405",
  1784 => x"0d747088",
  1785 => x"2a83fe80",
  1786 => x"06707298",
  1787 => x"2a077288",
  1788 => x"2b87fc80",
  1789 => x"80067398",
  1790 => x"2b81f00a",
  1791 => x"06717307",
  1792 => x"0780d5fc",
  1793 => x"0c565153",
  1794 => x"51028c05",
  1795 => x"0d0402f8",
  1796 => x"050d028e",
  1797 => x"0580f52d",
  1798 => x"74882b07",
  1799 => x"7083ffff",
  1800 => x"0680d5fc",
  1801 => x"0c510288",
  1802 => x"050d0402",
  1803 => x"ec050d76",
  1804 => x"787a5355",
  1805 => x"53815580",
  1806 => x"7125ae38",
  1807 => x"70527370",
  1808 => x"81055580",
  1809 => x"f52d7370",
  1810 => x"81055581",
  1811 => x"b72d7380",
  1812 => x"f52d5170",
  1813 => x"86387055",
  1814 => x"b8de0474",
  1815 => x"8638a073",
  1816 => x"81b72dff",
  1817 => x"125271d6",
  1818 => x"38807381",
  1819 => x"b72d0294",
  1820 => x"050d0402",
  1821 => x"e8050d77",
  1822 => x"56807056",
  1823 => x"54737624",
  1824 => x"b63880dd",
  1825 => x"8408742e",
  1826 => x"ae387351",
  1827 => x"b2862d80",
  1828 => x"d5fc0880",
  1829 => x"d5fc0809",
  1830 => x"81057080",
  1831 => x"d5fc0807",
  1832 => x"9f2a7705",
  1833 => x"81175757",
  1834 => x"53537476",
  1835 => x"24893880",
  1836 => x"dd840874",
  1837 => x"26d43872",
  1838 => x"80d5fc0c",
  1839 => x"0298050d",
  1840 => x"0402f005",
  1841 => x"0d80d5f8",
  1842 => x"081651b8",
  1843 => x"f32d80d5",
  1844 => x"fc08802e",
  1845 => x"9f388b53",
  1846 => x"80d5fc08",
  1847 => x"5280daf4",
  1848 => x"51b8ab2d",
  1849 => x"80ddb008",
  1850 => x"5473802e",
  1851 => x"873880da",
  1852 => x"f451732d",
  1853 => x"0290050d",
  1854 => x"0402dc05",
  1855 => x"0d80705a",
  1856 => x"557480d5",
  1857 => x"f80825b4",
  1858 => x"3880dd84",
  1859 => x"08752eac",
  1860 => x"387851b2",
  1861 => x"862d80d5",
  1862 => x"fc080981",
  1863 => x"057080d5",
  1864 => x"fc08079f",
  1865 => x"2a760581",
  1866 => x"1b5b5654",
  1867 => x"7480d5f8",
  1868 => x"08258938",
  1869 => x"80dd8408",
  1870 => x"7926d638",
  1871 => x"80557880",
  1872 => x"dd840827",
  1873 => x"81db3878",
  1874 => x"51b2862d",
  1875 => x"80d5fc08",
  1876 => x"802e81ad",
  1877 => x"3880d5fc",
  1878 => x"088b0580",
  1879 => x"f52d7084",
  1880 => x"2a708106",
  1881 => x"77107884",
  1882 => x"2b80daf4",
  1883 => x"0b80f52d",
  1884 => x"5c5c5351",
  1885 => x"55567380",
  1886 => x"2e80cb38",
  1887 => x"7416822b",
  1888 => x"bcc50b80",
  1889 => x"d4cc120c",
  1890 => x"54777531",
  1891 => x"1080ddb4",
  1892 => x"11555690",
  1893 => x"74708105",
  1894 => x"5681b72d",
  1895 => x"a07481b7",
  1896 => x"2d7681ff",
  1897 => x"06811658",
  1898 => x"5473802e",
  1899 => x"8a389c53",
  1900 => x"80daf452",
  1901 => x"bbbe048b",
  1902 => x"5380d5fc",
  1903 => x"085280dd",
  1904 => x"b61651bb",
  1905 => x"f9047416",
  1906 => x"822bb9c1",
  1907 => x"0b80d4cc",
  1908 => x"120c5476",
  1909 => x"81ff0681",
  1910 => x"16585473",
  1911 => x"802e8a38",
  1912 => x"9c5380da",
  1913 => x"f452bbf0",
  1914 => x"048b5380",
  1915 => x"d5fc0852",
  1916 => x"77753110",
  1917 => x"80ddb405",
  1918 => x"517655b8",
  1919 => x"ab2dbc96",
  1920 => x"04749029",
  1921 => x"75317010",
  1922 => x"80ddb405",
  1923 => x"515480d5",
  1924 => x"fc087481",
  1925 => x"b72d8119",
  1926 => x"59748b24",
  1927 => x"a338babe",
  1928 => x"04749029",
  1929 => x"75317010",
  1930 => x"80ddb405",
  1931 => x"8c773157",
  1932 => x"51548074",
  1933 => x"81b72d9e",
  1934 => x"14ff1656",
  1935 => x"5474f338",
  1936 => x"02a4050d",
  1937 => x"0402fc05",
  1938 => x"0d80d5f8",
  1939 => x"081351b8",
  1940 => x"f32d80d5",
  1941 => x"fc08802e",
  1942 => x"893880d5",
  1943 => x"fc0851a9",
  1944 => x"d32d800b",
  1945 => x"80d5f80c",
  1946 => x"b9f92d94",
  1947 => x"a52d0284",
  1948 => x"050d0402",
  1949 => x"f8050d73",
  1950 => x"5170fd2e",
  1951 => x"b13870fd",
  1952 => x"248a3870",
  1953 => x"fc2e80cd",
  1954 => x"38bdef04",
  1955 => x"70fe2eb8",
  1956 => x"3870ff2e",
  1957 => x"09810680",
  1958 => x"d63880d5",
  1959 => x"f8085170",
  1960 => x"802e80cb",
  1961 => x"38ff1180",
  1962 => x"d5f80cbd",
  1963 => x"ef0480d5",
  1964 => x"f808f405",
  1965 => x"7080d5f8",
  1966 => x"0c517080",
  1967 => x"25b13880",
  1968 => x"0b80d5f8",
  1969 => x"0cbdef04",
  1970 => x"80d5f808",
  1971 => x"810580d5",
  1972 => x"f80cbdef",
  1973 => x"0480d5f8",
  1974 => x"088c1170",
  1975 => x"80d5f80c",
  1976 => x"525280dd",
  1977 => x"84087126",
  1978 => x"86387180",
  1979 => x"d5f80cb9",
  1980 => x"f92d94a5",
  1981 => x"2d028805",
  1982 => x"0d0402fc",
  1983 => x"050d800b",
  1984 => x"80d5f80c",
  1985 => x"b9f92d93",
  1986 => x"882d80d5",
  1987 => x"fc0880d5",
  1988 => x"e80c80d4",
  1989 => x"c45195cb",
  1990 => x"2d028405",
  1991 => x"0d0402f8",
  1992 => x"050d810b",
  1993 => x"80ce8c0c",
  1994 => x"80d6a408",
  1995 => x"bff9ff06",
  1996 => x"81800770",
  1997 => x"80d6a40c",
  1998 => x"fc0c7351",
  1999 => x"bdfa2d02",
  2000 => x"88050d04",
  2001 => x"02f8050d",
  2002 => x"820b80ce",
  2003 => x"8c0c80d6",
  2004 => x"a408bffa",
  2005 => x"ff068280",
  2006 => x"077080d6",
  2007 => x"a40cfc0c",
  2008 => x"7351bdfa",
  2009 => x"2d028805",
  2010 => x"0d0402f8",
  2011 => x"050d830b",
  2012 => x"80ce8c0c",
  2013 => x"80d6a408",
  2014 => x"bfffff06",
  2015 => x"87800770",
  2016 => x"80d6a40c",
  2017 => x"fc0c7351",
  2018 => x"bdfa2d02",
  2019 => x"88050d04",
  2020 => x"7180ddb0",
  2021 => x"0c040000",
  2022 => x"00ffffff",
  2023 => x"ff00ffff",
  2024 => x"ffff00ff",
  2025 => x"ffffff00",
  2026 => x"54686572",
  2027 => x"65206973",
  2028 => x"206e6f20",
  2029 => x"696d6167",
  2030 => x"65207768",
  2031 => x"656e206c",
  2032 => x"6f616469",
  2033 => x"6e670000",
  2034 => x"436f6e74",
  2035 => x"696e7565",
  2036 => x"00000000",
  2037 => x"3d205a58",
  2038 => x"38312f5a",
  2039 => x"58383020",
  2040 => x"436f6e66",
  2041 => x"69677572",
  2042 => x"6174696f",
  2043 => x"6e203d00",
  2044 => x"3d3d3d3d",
  2045 => x"3d3d3d3d",
  2046 => x"3d3d3d3d",
  2047 => x"3d3d3d3d",
  2048 => x"3d3d3d3d",
  2049 => x"3d3d3d3d",
  2050 => x"3d3d3d00",
  2051 => x"4c6f7720",
  2052 => x"52414d3a",
  2053 => x"204f6666",
  2054 => x"2f384b42",
  2055 => x"00000000",
  2056 => x"51532043",
  2057 => x"4852533a",
  2058 => x"44697361",
  2059 => x"626c6564",
  2060 => x"2f456e61",
  2061 => x"626c6564",
  2062 => x"28463129",
  2063 => x"00000000",
  2064 => x"4348524f",
  2065 => x"4d413831",
  2066 => x"3a204469",
  2067 => x"7361626c",
  2068 => x"65642f45",
  2069 => x"6e61626c",
  2070 => x"65640000",
  2071 => x"496e7665",
  2072 => x"72736520",
  2073 => x"76696465",
  2074 => x"6f3a204f",
  2075 => x"66662f4f",
  2076 => x"6e000000",
  2077 => x"426c6163",
  2078 => x"6b20626f",
  2079 => x"72646572",
  2080 => x"3a204f66",
  2081 => x"662f4f6e",
  2082 => x"00000000",
  2083 => x"56696465",
  2084 => x"6f206672",
  2085 => x"65717565",
  2086 => x"6e63793a",
  2087 => x"20353048",
  2088 => x"7a2f3630",
  2089 => x"487a0000",
  2090 => x"476f2042",
  2091 => x"61636b00",
  2092 => x"536c6f77",
  2093 => x"206d6f64",
  2094 => x"65207370",
  2095 => x"6565643a",
  2096 => x"204f7269",
  2097 => x"67696e61",
  2098 => x"6c000000",
  2099 => x"536c6f77",
  2100 => x"206d6f64",
  2101 => x"65207370",
  2102 => x"6565643a",
  2103 => x"204e6f57",
  2104 => x"61697400",
  2105 => x"536c6f77",
  2106 => x"206d6f64",
  2107 => x"65207370",
  2108 => x"6565643a",
  2109 => x"20783200",
  2110 => x"536c6f77",
  2111 => x"206d6f64",
  2112 => x"65207370",
  2113 => x"6565643a",
  2114 => x"20783800",
  2115 => x"43485224",
  2116 => x"3132382f",
  2117 => x"5544473a",
  2118 => x"20313238",
  2119 => x"20436861",
  2120 => x"72730000",
  2121 => x"43485224",
  2122 => x"3132382f",
  2123 => x"5544473a",
  2124 => x"20363420",
  2125 => x"43686172",
  2126 => x"73000000",
  2127 => x"43485224",
  2128 => x"3132382f",
  2129 => x"5544473a",
  2130 => x"20446973",
  2131 => x"61626c65",
  2132 => x"64000000",
  2133 => x"4a6f7973",
  2134 => x"7469636b",
  2135 => x"3a204375",
  2136 => x"72736f72",
  2137 => x"00000000",
  2138 => x"4a6f7973",
  2139 => x"7469636b",
  2140 => x"3a205369",
  2141 => x"6e636c61",
  2142 => x"69720000",
  2143 => x"4a6f7973",
  2144 => x"7469636b",
  2145 => x"3a205a58",
  2146 => x"38310000",
  2147 => x"4d61696e",
  2148 => x"2052414d",
  2149 => x"3a203136",
  2150 => x"4b420000",
  2151 => x"4d61696e",
  2152 => x"2052414d",
  2153 => x"3a203332",
  2154 => x"4b420000",
  2155 => x"4d61696e",
  2156 => x"2052414d",
  2157 => x"3a203438",
  2158 => x"4b420000",
  2159 => x"4d61696e",
  2160 => x"2052414d",
  2161 => x"3a20314b",
  2162 => x"42000000",
  2163 => x"436f6d70",
  2164 => x"75746572",
  2165 => x"204d6f64",
  2166 => x"656c3a20",
  2167 => x"5a583831",
  2168 => x"00000000",
  2169 => x"436f6d70",
  2170 => x"75746572",
  2171 => x"204d6f64",
  2172 => x"656c3a20",
  2173 => x"5a583830",
  2174 => x"00000000",
  2175 => x"3d3d205a",
  2176 => x"5838312f",
  2177 => x"5a583830",
  2178 => x"20666f72",
  2179 => x"205a5844",
  2180 => x"4f53203d",
  2181 => x"3d000000",
  2182 => x"3d3d3d3d",
  2183 => x"3d3d3d3d",
  2184 => x"3d3d3d3d",
  2185 => x"3d3d3d3d",
  2186 => x"3d3d3d3d",
  2187 => x"3d3d3d3d",
  2188 => x"3d000000",
  2189 => x"52657365",
  2190 => x"74000000",
  2191 => x"4c6f6164",
  2192 => x"20546170",
  2193 => x"6520282e",
  2194 => x"70292010",
  2195 => x"00000000",
  2196 => x"4c6f6164",
  2197 => x"20546170",
  2198 => x"6520282e",
  2199 => x"6f292010",
  2200 => x"00000000",
  2201 => x"4c6f6164",
  2202 => x"20526f6d",
  2203 => x"2020282e",
  2204 => x"726f6d29",
  2205 => x"20100000",
  2206 => x"436f6e66",
  2207 => x"69677572",
  2208 => x"6174696f",
  2209 => x"6e206f70",
  2210 => x"74696f6e",
  2211 => x"73201000",
  2212 => x"4b657962",
  2213 => x"6f617264",
  2214 => x"2048656c",
  2215 => x"70000000",
  2216 => x"45786974",
  2217 => x"00000000",
  2218 => x"3d3d205a",
  2219 => x"5838312f",
  2220 => x"5a583830",
  2221 => x"20666f72",
  2222 => x"205a5855",
  2223 => x"4e4f203d",
  2224 => x"3d000000",
  2225 => x"524f4d20",
  2226 => x"6c6f6164",
  2227 => x"696e6720",
  2228 => x"6661696c",
  2229 => x"65640000",
  2230 => x"4f4b0000",
  2231 => x"54617065",
  2232 => x"2066696c",
  2233 => x"65204c6f",
  2234 => x"61646564",
  2235 => x"2e000000",
  2236 => x"54797065",
  2237 => x"204c4f41",
  2238 => x"44202222",
  2239 => x"202b2045",
  2240 => x"4e544552",
  2241 => x"206f6e20",
  2242 => x"5a583831",
  2243 => x"00000000",
  2244 => x"3d205a58",
  2245 => x"38312f5a",
  2246 => x"58383020",
  2247 => x"4b657962",
  2248 => x"6f617264",
  2249 => x"2048656c",
  2250 => x"70203d00",
  2251 => x"5363726f",
  2252 => x"6c6c204c",
  2253 => x"6f636b3a",
  2254 => x"20636861",
  2255 => x"6e676520",
  2256 => x"62657477",
  2257 => x"65656e00",
  2258 => x"52474220",
  2259 => x"616e6420",
  2260 => x"56474120",
  2261 => x"76696465",
  2262 => x"6f206d6f",
  2263 => x"64650000",
  2264 => x"4374726c",
  2265 => x"2b416c74",
  2266 => x"2b44656c",
  2267 => x"6574653a",
  2268 => x"20536f66",
  2269 => x"74205265",
  2270 => x"73657400",
  2271 => x"4374726c",
  2272 => x"2b416c74",
  2273 => x"2b426163",
  2274 => x"6b737061",
  2275 => x"63653a20",
  2276 => x"48617264",
  2277 => x"20726573",
  2278 => x"65740000",
  2279 => x"45736320",
  2280 => x"6f72206a",
  2281 => x"6f797374",
  2282 => x"69636b20",
  2283 => x"62742e32",
  2284 => x"3a20746f",
  2285 => x"2073686f",
  2286 => x"77000000",
  2287 => x"6f722068",
  2288 => x"69646520",
  2289 => x"74686520",
  2290 => x"6f707469",
  2291 => x"6f6e7320",
  2292 => x"6d656e75",
  2293 => x"2e000000",
  2294 => x"57415344",
  2295 => x"202f2063",
  2296 => x"7572736f",
  2297 => x"72206b65",
  2298 => x"7973202f",
  2299 => x"206a6f79",
  2300 => x"73746963",
  2301 => x"6b000000",
  2302 => x"746f2073",
  2303 => x"656c6563",
  2304 => x"74206d65",
  2305 => x"6e75206f",
  2306 => x"7074696f",
  2307 => x"6e2e0000",
  2308 => x"456e7465",
  2309 => x"72202f20",
  2310 => x"46697265",
  2311 => x"20746f20",
  2312 => x"63686f6f",
  2313 => x"7365206f",
  2314 => x"7074696f",
  2315 => x"6e2e0000",
  2316 => x"3d205a58",
  2317 => x"38312f5a",
  2318 => x"58383020",
  2319 => x"436f7265",
  2320 => x"20437265",
  2321 => x"64697473",
  2322 => x"20203d00",
  2323 => x"5a583831",
  2324 => x"2f5a5838",
  2325 => x"3020636f",
  2326 => x"72652066",
  2327 => x"6f72205a",
  2328 => x"58554e4f",
  2329 => x"2c200000",
  2330 => x"5a58444f",
  2331 => x"5320616e",
  2332 => x"64205a58",
  2333 => x"444f532b",
  2334 => x"20626f61",
  2335 => x"7264732e",
  2336 => x"00000000",
  2337 => x"4f726967",
  2338 => x"696e616c",
  2339 => x"20636f72",
  2340 => x"65732062",
  2341 => x"793a0000",
  2342 => x"202d2053",
  2343 => x"7a6f6d62",
  2344 => x"61746865",
  2345 => x"6c796920",
  2346 => x"47796f72",
  2347 => x"67792028",
  2348 => x"4d697374",
  2349 => x"29000000",
  2350 => x"202d2053",
  2351 => x"6f726765",
  2352 => x"6c696720",
  2353 => x"284d6973",
  2354 => x"74657229",
  2355 => x"00000000",
  2356 => x"506f7274",
  2357 => x"206d6164",
  2358 => x"65206279",
  2359 => x"3a204176",
  2360 => x"6c697841",
  2361 => x"00000000",
  2362 => x"496e6974",
  2363 => x"69616c69",
  2364 => x"7a696e67",
  2365 => x"20534420",
  2366 => x"63617264",
  2367 => x"0a000000",
  2368 => x"4c6f6164",
  2369 => x"696e6720",
  2370 => x"696e6974",
  2371 => x"69616c20",
  2372 => x"524f4d2e",
  2373 => x"2e2e0a00",
  2374 => x"5a583831",
  2375 => x"20202020",
  2376 => x"20202000",
  2377 => x"524f4d53",
  2378 => x"20202020",
  2379 => x"20202000",
  2380 => x"5a583858",
  2381 => x"20202020",
  2382 => x"524f4d00",
  2383 => x"4572726f",
  2384 => x"72204c6f",
  2385 => x"6164696e",
  2386 => x"6720524f",
  2387 => x"4d2e2e2e",
  2388 => x"0a000000",
  2389 => x"2e2e2020",
  2390 => x"20202020",
  2391 => x"20202000",
  2392 => x"16200000",
  2393 => x"14200000",
  2394 => x"15200000",
  2395 => x"53442069",
  2396 => x"6e69742e",
  2397 => x"2e2e0a00",
  2398 => x"53442063",
  2399 => x"61726420",
  2400 => x"72657365",
  2401 => x"74206661",
  2402 => x"696c6564",
  2403 => x"210a0000",
  2404 => x"53444843",
  2405 => x"20657272",
  2406 => x"6f72210a",
  2407 => x"00000000",
  2408 => x"57726974",
  2409 => x"65206661",
  2410 => x"696c6564",
  2411 => x"0a000000",
  2412 => x"52656164",
  2413 => x"20666169",
  2414 => x"6c65640a",
  2415 => x"00000000",
  2416 => x"43617264",
  2417 => x"20696e69",
  2418 => x"74206661",
  2419 => x"696c6564",
  2420 => x"0a000000",
  2421 => x"46415431",
  2422 => x"36202020",
  2423 => x"00000000",
  2424 => x"46415433",
  2425 => x"32202020",
  2426 => x"00000000",
  2427 => x"4e6f2070",
  2428 => x"61727469",
  2429 => x"74696f6e",
  2430 => x"20736967",
  2431 => x"0a000000",
  2432 => x"42616420",
  2433 => x"70617274",
  2434 => x"0a000000",
  2435 => x"4261636b",
  2436 => x"00000000",
  2437 => x"00000002",
  2438 => x"00000002",
  2439 => x"00001fd4",
  2440 => x"00000342",
  2441 => x"00000002",
  2442 => x"00001ff0",
  2443 => x"00000342",
  2444 => x"00000003",
  2445 => x"00002704",
  2446 => x"00000002",
  2447 => x"00000003",
  2448 => x"000026f4",
  2449 => x"00000004",
  2450 => x"00000001",
  2451 => x"0000200c",
  2452 => x"00000000",
  2453 => x"00000003",
  2454 => x"000026e8",
  2455 => x"00000003",
  2456 => x"00000001",
  2457 => x"00002020",
  2458 => x"00000001",
  2459 => x"00000003",
  2460 => x"000026dc",
  2461 => x"00000003",
  2462 => x"00000001",
  2463 => x"00002040",
  2464 => x"00000002",
  2465 => x"00000001",
  2466 => x"0000205c",
  2467 => x"00000003",
  2468 => x"00000001",
  2469 => x"00002074",
  2470 => x"00000004",
  2471 => x"00000003",
  2472 => x"000026cc",
  2473 => x"00000003",
  2474 => x"00000001",
  2475 => x"0000208c",
  2476 => x"00000005",
  2477 => x"00000004",
  2478 => x"000020a8",
  2479 => x"00002b28",
  2480 => x"00000000",
  2481 => x"00000000",
  2482 => x"00000000",
  2483 => x"000020b0",
  2484 => x"000020cc",
  2485 => x"000020e4",
  2486 => x"000020f8",
  2487 => x"0000210c",
  2488 => x"00002124",
  2489 => x"0000213c",
  2490 => x"00002154",
  2491 => x"00002168",
  2492 => x"0000217c",
  2493 => x"0000218c",
  2494 => x"0000219c",
  2495 => x"000021ac",
  2496 => x"000021bc",
  2497 => x"000021cc",
  2498 => x"000021e4",
  2499 => x"00000000",
  2500 => x"00000002",
  2501 => x"000021fc",
  2502 => x"00000343",
  2503 => x"00000002",
  2504 => x"00002218",
  2505 => x"00000343",
  2506 => x"00000002",
  2507 => x"00002234",
  2508 => x"00000386",
  2509 => x"00000002",
  2510 => x"0000223c",
  2511 => x"00001f1e",
  2512 => x"00000002",
  2513 => x"00002250",
  2514 => x"00001f44",
  2515 => x"00000002",
  2516 => x"00002264",
  2517 => x"00001f6a",
  2518 => x"00000002",
  2519 => x"00002278",
  2520 => x"00000353",
  2521 => x"00000002",
  2522 => x"00002290",
  2523 => x"00000363",
  2524 => x"00000002",
  2525 => x"000022a0",
  2526 => x"000009a5",
  2527 => x"00000000",
  2528 => x"00000000",
  2529 => x"00000000",
  2530 => x"00000002",
  2531 => x"000022a8",
  2532 => x"00000343",
  2533 => x"00000002",
  2534 => x"00002218",
  2535 => x"00000343",
  2536 => x"00000002",
  2537 => x"00002234",
  2538 => x"00000386",
  2539 => x"00000002",
  2540 => x"0000223c",
  2541 => x"00001f1e",
  2542 => x"00000002",
  2543 => x"00002250",
  2544 => x"00001f44",
  2545 => x"00000002",
  2546 => x"00002264",
  2547 => x"00001f6a",
  2548 => x"00000002",
  2549 => x"00002278",
  2550 => x"00000353",
  2551 => x"00000002",
  2552 => x"00002290",
  2553 => x"00000363",
  2554 => x"00000002",
  2555 => x"000022a0",
  2556 => x"000009a5",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000000",
  2560 => x"00000004",
  2561 => x"000022c4",
  2562 => x"00002800",
  2563 => x"00000004",
  2564 => x"000022d8",
  2565 => x"00002b28",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000004",
  2570 => x"000022dc",
  2571 => x"00002824",
  2572 => x"00000004",
  2573 => x"000022f0",
  2574 => x"00002824",
  2575 => x"00000004",
  2576 => x"0000259c",
  2577 => x"00002824",
  2578 => x"00000004",
  2579 => x"00001fa8",
  2580 => x"00002824",
  2581 => x"00000004",
  2582 => x"0000259c",
  2583 => x"00002824",
  2584 => x"00000004",
  2585 => x"00001fc8",
  2586 => x"00002b28",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000002",
  2591 => x"00002310",
  2592 => x"00000342",
  2593 => x"00000002",
  2594 => x"00001ff0",
  2595 => x"00000342",
  2596 => x"00000002",
  2597 => x"0000232c",
  2598 => x"00000342",
  2599 => x"00000002",
  2600 => x"00002348",
  2601 => x"00000342",
  2602 => x"00000002",
  2603 => x"00002360",
  2604 => x"00000342",
  2605 => x"00000002",
  2606 => x"0000237c",
  2607 => x"00000342",
  2608 => x"00000002",
  2609 => x"0000239c",
  2610 => x"00000342",
  2611 => x"00000002",
  2612 => x"000023bc",
  2613 => x"00000342",
  2614 => x"00000002",
  2615 => x"000023d8",
  2616 => x"00000342",
  2617 => x"00000002",
  2618 => x"000023f8",
  2619 => x"00000342",
  2620 => x"00000002",
  2621 => x"00002410",
  2622 => x"00000342",
  2623 => x"00000002",
  2624 => x"0000259c",
  2625 => x"00000342",
  2626 => x"00000004",
  2627 => x"000022d8",
  2628 => x"00002b28",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000002",
  2633 => x"00002430",
  2634 => x"00000342",
  2635 => x"00000002",
  2636 => x"00001ff0",
  2637 => x"00000342",
  2638 => x"00000002",
  2639 => x"0000244c",
  2640 => x"00000342",
  2641 => x"00000002",
  2642 => x"00002468",
  2643 => x"00000342",
  2644 => x"00000002",
  2645 => x"0000259c",
  2646 => x"00000342",
  2647 => x"00000002",
  2648 => x"00002484",
  2649 => x"00000342",
  2650 => x"00000002",
  2651 => x"00002498",
  2652 => x"00000342",
  2653 => x"00000002",
  2654 => x"000024b8",
  2655 => x"00000342",
  2656 => x"00000002",
  2657 => x"0000259c",
  2658 => x"00000342",
  2659 => x"00000002",
  2660 => x"000024d0",
  2661 => x"00000342",
  2662 => x"00000002",
  2663 => x"0000259c",
  2664 => x"00000342",
  2665 => x"00000002",
  2666 => x"0000259c",
  2667 => x"00000342",
  2668 => x"00000004",
  2669 => x"000022d8",
  2670 => x"00002b28",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000006",
  2693 => x"00000043",
  2694 => x"00000042",
  2695 => x"0000003b",
  2696 => x"0000004b",
  2697 => x"0000007e",
  2698 => x"00000003",
  2699 => x"0000000b",
  2700 => x"00000083",
  2701 => x"00000023",
  2702 => x"0000007e",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000002",
  2706 => x"00002eb4",
  2707 => x"00001cc1",
  2708 => x"00000002",
  2709 => x"00002ed2",
  2710 => x"00001cc1",
  2711 => x"00000002",
  2712 => x"00002ef0",
  2713 => x"00001cc1",
  2714 => x"00000002",
  2715 => x"00002f0e",
  2716 => x"00001cc1",
  2717 => x"00000002",
  2718 => x"00002f2c",
  2719 => x"00001cc1",
  2720 => x"00000002",
  2721 => x"00002f4a",
  2722 => x"00001cc1",
  2723 => x"00000002",
  2724 => x"00002f68",
  2725 => x"00001cc1",
  2726 => x"00000002",
  2727 => x"00002f86",
  2728 => x"00001cc1",
  2729 => x"00000002",
  2730 => x"00002fa4",
  2731 => x"00001cc1",
  2732 => x"00000002",
  2733 => x"00002fc2",
  2734 => x"00001cc1",
  2735 => x"00000002",
  2736 => x"00002fe0",
  2737 => x"00001cc1",
  2738 => x"00000002",
  2739 => x"00002ffe",
  2740 => x"00001cc1",
  2741 => x"00000002",
  2742 => x"0000301c",
  2743 => x"00001cc1",
  2744 => x"00000004",
  2745 => x"0000260c",
  2746 => x"00000000",
  2747 => x"00000000",
  2748 => x"00000000",
  2749 => x"00001e73",
  2750 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

